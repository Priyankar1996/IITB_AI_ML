-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_34_start: Boolean;
  signal convTranspose_CP_34_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_ConvTranspose_input_pipe_746_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1090_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_746_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_746_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_993_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1084_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_978_inst_req_1 : boolean;
  signal type_cast_732_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_746_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_993_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_593_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1063_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1016_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1016_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_593_inst_req_1 : boolean;
  signal type_cast_732_inst_ack_0 : boolean;
  signal addr_of_694_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_req_1 : boolean;
  signal ptr_deref_623_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_ack_1 : boolean;
  signal type_cast_597_inst_ack_1 : boolean;
  signal type_cast_597_inst_req_1 : boolean;
  signal type_cast_597_inst_req_0 : boolean;
  signal type_cast_597_inst_ack_0 : boolean;
  signal type_cast_543_inst_ack_1 : boolean;
  signal type_cast_543_inst_req_1 : boolean;
  signal type_cast_543_inst_ack_0 : boolean;
  signal type_cast_543_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1056_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_40_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1019_inst_req_1 : boolean;
  signal addr_of_694_final_reg_req_1 : boolean;
  signal type_cast_44_inst_req_0 : boolean;
  signal type_cast_44_inst_ack_0 : boolean;
  signal type_cast_44_inst_req_1 : boolean;
  signal type_cast_44_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_987_inst_ack_1 : boolean;
  signal type_cast_1396_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1075_inst_req_0 : boolean;
  signal type_cast_144_inst_req_0 : boolean;
  signal type_cast_144_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1002_inst_req_1 : boolean;
  signal if_stmt_637_branch_req_0 : boolean;
  signal WPIPE_Block1_start_1019_inst_ack_1 : boolean;
  signal type_cast_57_inst_req_0 : boolean;
  signal type_cast_57_inst_ack_0 : boolean;
  signal type_cast_57_inst_req_1 : boolean;
  signal ptr_deref_623_store_0_req_1 : boolean;
  signal type_cast_57_inst_ack_1 : boolean;
  signal type_cast_1396_inst_req_1 : boolean;
  signal type_cast_1426_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_65_inst_req_0 : boolean;
  signal WPIPE_Block0_start_996_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_65_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_593_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_65_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_65_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1069_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1022_inst_req_0 : boolean;
  signal type_cast_615_inst_ack_1 : boolean;
  signal type_cast_69_inst_req_0 : boolean;
  signal type_cast_69_inst_ack_0 : boolean;
  signal type_cast_69_inst_req_1 : boolean;
  signal type_cast_69_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_593_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1063_inst_req_1 : boolean;
  signal type_cast_1426_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_78_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_728_inst_ack_1 : boolean;
  signal type_cast_615_inst_req_1 : boolean;
  signal type_cast_82_inst_req_0 : boolean;
  signal WPIPE_Block0_start_978_inst_ack_1 : boolean;
  signal type_cast_82_inst_ack_0 : boolean;
  signal array_obj_ref_693_index_offset_ack_1 : boolean;
  signal type_cast_82_inst_req_1 : boolean;
  signal type_cast_82_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1063_inst_ack_0 : boolean;
  signal type_cast_664_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_978_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_90_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_90_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_90_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_90_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_710_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_710_inst_req_1 : boolean;
  signal addr_of_694_final_reg_ack_0 : boolean;
  signal type_cast_714_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1022_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1037_inst_req_0 : boolean;
  signal type_cast_94_inst_req_0 : boolean;
  signal type_cast_94_inst_ack_0 : boolean;
  signal array_obj_ref_693_index_offset_req_1 : boolean;
  signal type_cast_94_inst_req_1 : boolean;
  signal ptr_deref_623_store_0_ack_0 : boolean;
  signal type_cast_94_inst_ack_1 : boolean;
  signal type_cast_664_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_697_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_req_1 : boolean;
  signal ptr_deref_623_store_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_103_inst_ack_1 : boolean;
  signal type_cast_1436_inst_ack_0 : boolean;
  signal type_cast_714_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1063_inst_ack_1 : boolean;
  signal type_cast_107_inst_req_0 : boolean;
  signal type_cast_107_inst_ack_0 : boolean;
  signal type_cast_107_inst_req_1 : boolean;
  signal type_cast_107_inst_ack_1 : boolean;
  signal type_cast_664_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_697_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_115_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_115_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_115_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_115_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_728_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_710_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_710_inst_req_0 : boolean;
  signal addr_of_694_final_reg_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1301_inst_ack_0 : boolean;
  signal type_cast_615_inst_ack_0 : boolean;
  signal type_cast_119_inst_req_0 : boolean;
  signal type_cast_119_inst_ack_0 : boolean;
  signal type_cast_119_inst_req_1 : boolean;
  signal type_cast_119_inst_ack_1 : boolean;
  signal type_cast_732_inst_ack_1 : boolean;
  signal type_cast_664_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_ack_0 : boolean;
  signal type_cast_579_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_128_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1069_inst_ack_1 : boolean;
  signal type_cast_615_inst_req_0 : boolean;
  signal array_obj_ref_693_index_offset_ack_0 : boolean;
  signal type_cast_132_inst_req_0 : boolean;
  signal type_cast_132_inst_ack_0 : boolean;
  signal array_obj_ref_693_index_offset_req_0 : boolean;
  signal type_cast_132_inst_req_1 : boolean;
  signal type_cast_132_inst_ack_1 : boolean;
  signal type_cast_732_inst_req_1 : boolean;
  signal type_cast_579_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_697_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_ack_1 : boolean;
  signal type_cast_345_inst_req_1 : boolean;
  signal type_cast_345_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_981_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1025_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_354_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_354_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_354_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_354_inst_ack_1 : boolean;
  signal type_cast_358_inst_req_0 : boolean;
  signal type_cast_144_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_539_inst_ack_1 : boolean;
  signal type_cast_144_inst_ack_1 : boolean;
  signal type_cast_714_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_697_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_ack_0 : boolean;
  signal type_cast_579_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1056_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_153_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_987_inst_req_1 : boolean;
  signal type_cast_157_inst_req_0 : boolean;
  signal type_cast_157_inst_ack_0 : boolean;
  signal type_cast_157_inst_req_1 : boolean;
  signal type_cast_157_inst_ack_1 : boolean;
  signal type_cast_714_inst_req_1 : boolean;
  signal type_cast_579_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_165_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_165_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_165_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_165_inst_ack_1 : boolean;
  signal type_cast_169_inst_req_0 : boolean;
  signal type_cast_169_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1019_inst_req_0 : boolean;
  signal type_cast_169_inst_req_1 : boolean;
  signal type_cast_169_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_178_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_978_inst_req_0 : boolean;
  signal type_cast_182_inst_req_0 : boolean;
  signal type_cast_182_inst_ack_0 : boolean;
  signal type_cast_182_inst_req_1 : boolean;
  signal type_cast_182_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_539_inst_req_1 : boolean;
  signal if_stmt_637_branch_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_190_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_728_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1022_inst_req_1 : boolean;
  signal type_cast_194_inst_req_0 : boolean;
  signal type_cast_194_inst_ack_0 : boolean;
  signal type_cast_194_inst_req_1 : boolean;
  signal type_cast_194_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_575_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_575_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1002_inst_ack_1 : boolean;
  signal type_cast_701_inst_ack_1 : boolean;
  signal type_cast_207_inst_req_0 : boolean;
  signal type_cast_207_inst_ack_0 : boolean;
  signal type_cast_207_inst_req_1 : boolean;
  signal type_cast_207_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1022_inst_ack_1 : boolean;
  signal type_cast_216_inst_req_0 : boolean;
  signal type_cast_216_inst_ack_0 : boolean;
  signal type_cast_216_inst_req_1 : boolean;
  signal type_cast_216_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_575_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_575_inst_req_0 : boolean;
  signal WPIPE_Block0_start_996_inst_req_1 : boolean;
  signal type_cast_220_inst_req_0 : boolean;
  signal type_cast_220_inst_ack_0 : boolean;
  signal type_cast_220_inst_req_1 : boolean;
  signal type_cast_220_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_611_inst_ack_1 : boolean;
  signal type_cast_224_inst_req_0 : boolean;
  signal type_cast_224_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_539_inst_ack_0 : boolean;
  signal type_cast_224_inst_req_1 : boolean;
  signal type_cast_224_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_611_inst_req_1 : boolean;
  signal type_cast_261_inst_req_0 : boolean;
  signal type_cast_261_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_539_inst_req_0 : boolean;
  signal type_cast_261_inst_req_1 : boolean;
  signal type_cast_261_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1006_inst_req_1 : boolean;
  signal type_cast_1396_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_611_inst_ack_0 : boolean;
  signal type_cast_265_inst_req_0 : boolean;
  signal type_cast_265_inst_ack_0 : boolean;
  signal type_cast_265_inst_req_1 : boolean;
  signal type_cast_265_inst_ack_1 : boolean;
  signal type_cast_561_inst_ack_1 : boolean;
  signal type_cast_561_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_611_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1056_inst_req_1 : boolean;
  signal type_cast_269_inst_req_0 : boolean;
  signal type_cast_269_inst_ack_0 : boolean;
  signal type_cast_269_inst_req_1 : boolean;
  signal type_cast_269_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1301_inst_req_0 : boolean;
  signal type_cast_273_inst_req_0 : boolean;
  signal type_cast_273_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1019_inst_ack_0 : boolean;
  signal type_cast_273_inst_req_1 : boolean;
  signal type_cast_273_inst_ack_1 : boolean;
  signal type_cast_561_inst_ack_0 : boolean;
  signal type_cast_561_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_291_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_728_inst_req_0 : boolean;
  signal type_cast_701_inst_req_1 : boolean;
  signal type_cast_295_inst_req_0 : boolean;
  signal type_cast_295_inst_ack_0 : boolean;
  signal type_cast_295_inst_req_1 : boolean;
  signal type_cast_295_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_304_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_304_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_304_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_304_inst_ack_1 : boolean;
  signal type_cast_701_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1034_inst_req_1 : boolean;
  signal type_cast_308_inst_req_0 : boolean;
  signal type_cast_308_inst_ack_0 : boolean;
  signal type_cast_308_inst_req_1 : boolean;
  signal type_cast_308_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_557_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_996_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_557_inst_req_1 : boolean;
  signal if_stmt_637_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_316_inst_ack_1 : boolean;
  signal type_cast_701_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1034_inst_ack_1 : boolean;
  signal type_cast_320_inst_req_0 : boolean;
  signal type_cast_320_inst_ack_0 : boolean;
  signal type_cast_320_inst_req_1 : boolean;
  signal type_cast_320_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_557_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_329_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1056_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_329_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_557_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_329_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_329_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1025_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1025_inst_ack_0 : boolean;
  signal type_cast_333_inst_req_0 : boolean;
  signal type_cast_333_inst_ack_0 : boolean;
  signal type_cast_333_inst_req_1 : boolean;
  signal type_cast_333_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_996_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_341_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_341_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_341_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_341_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1025_inst_req_1 : boolean;
  signal type_cast_345_inst_req_0 : boolean;
  signal type_cast_345_inst_ack_0 : boolean;
  signal type_cast_358_inst_ack_0 : boolean;
  signal type_cast_358_inst_req_1 : boolean;
  signal type_cast_358_inst_ack_1 : boolean;
  signal ptr_deref_1372_load_0_ack_1 : boolean;
  signal WPIPE_Block0_start_981_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_366_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_990_inst_req_0 : boolean;
  signal type_cast_370_inst_req_0 : boolean;
  signal type_cast_370_inst_ack_0 : boolean;
  signal type_cast_370_inst_req_1 : boolean;
  signal type_cast_370_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_379_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_379_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_379_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_379_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_990_inst_ack_0 : boolean;
  signal type_cast_383_inst_req_0 : boolean;
  signal type_cast_383_inst_ack_0 : boolean;
  signal type_cast_383_inst_req_1 : boolean;
  signal type_cast_383_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_981_inst_req_1 : boolean;
  signal WPIPE_Block0_start_981_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_391_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_391_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_391_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_391_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_999_inst_req_0 : boolean;
  signal WPIPE_Block0_start_999_inst_ack_0 : boolean;
  signal type_cast_395_inst_req_0 : boolean;
  signal type_cast_395_inst_ack_0 : boolean;
  signal type_cast_395_inst_req_1 : boolean;
  signal type_cast_395_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1028_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_404_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_404_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_404_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_404_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1028_inst_ack_0 : boolean;
  signal type_cast_408_inst_req_0 : boolean;
  signal type_cast_408_inst_ack_0 : boolean;
  signal type_cast_408_inst_req_1 : boolean;
  signal type_cast_408_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1006_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1006_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_999_inst_req_1 : boolean;
  signal WPIPE_Block0_start_999_inst_ack_1 : boolean;
  signal if_stmt_421_branch_req_0 : boolean;
  signal if_stmt_421_branch_ack_1 : boolean;
  signal if_stmt_421_branch_ack_0 : boolean;
  signal if_stmt_436_branch_req_0 : boolean;
  signal if_stmt_436_branch_ack_1 : boolean;
  signal if_stmt_436_branch_ack_0 : boolean;
  signal type_cast_457_inst_req_0 : boolean;
  signal type_cast_457_inst_ack_0 : boolean;
  signal type_cast_457_inst_req_1 : boolean;
  signal type_cast_457_inst_ack_1 : boolean;
  signal array_obj_ref_486_index_offset_req_0 : boolean;
  signal array_obj_ref_486_index_offset_ack_0 : boolean;
  signal array_obj_ref_486_index_offset_req_1 : boolean;
  signal array_obj_ref_486_index_offset_ack_1 : boolean;
  signal addr_of_487_final_reg_req_0 : boolean;
  signal addr_of_487_final_reg_ack_0 : boolean;
  signal addr_of_487_final_reg_req_1 : boolean;
  signal addr_of_487_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_490_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_490_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_490_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_490_inst_ack_1 : boolean;
  signal type_cast_494_inst_req_0 : boolean;
  signal type_cast_494_inst_ack_0 : boolean;
  signal type_cast_494_inst_req_1 : boolean;
  signal type_cast_494_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_503_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_503_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_503_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_503_inst_ack_1 : boolean;
  signal type_cast_507_inst_req_0 : boolean;
  signal type_cast_507_inst_ack_0 : boolean;
  signal type_cast_507_inst_req_1 : boolean;
  signal type_cast_507_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_521_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_521_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_521_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_521_inst_ack_1 : boolean;
  signal type_cast_525_inst_req_0 : boolean;
  signal type_cast_525_inst_ack_0 : boolean;
  signal type_cast_525_inst_req_1 : boolean;
  signal type_cast_525_inst_ack_1 : boolean;
  signal type_cast_750_inst_req_0 : boolean;
  signal type_cast_750_inst_ack_0 : boolean;
  signal type_cast_750_inst_req_1 : boolean;
  signal type_cast_750_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1093_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_764_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_764_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_764_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_764_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1090_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1084_inst_req_1 : boolean;
  signal type_cast_1338_inst_ack_1 : boolean;
  signal type_cast_768_inst_req_0 : boolean;
  signal type_cast_768_inst_ack_0 : boolean;
  signal type_cast_768_inst_req_1 : boolean;
  signal type_cast_768_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_993_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1066_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_782_inst_req_0 : boolean;
  signal type_cast_1054_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_782_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_993_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_782_inst_req_1 : boolean;
  signal type_cast_1054_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_782_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1090_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1084_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1016_inst_ack_0 : boolean;
  signal type_cast_1396_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1016_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1286_inst_ack_1 : boolean;
  signal type_cast_786_inst_req_0 : boolean;
  signal type_cast_786_inst_ack_0 : boolean;
  signal type_cast_786_inst_req_1 : boolean;
  signal type_cast_786_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1066_inst_req_1 : boolean;
  signal type_cast_1426_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_800_inst_req_0 : boolean;
  signal type_cast_1054_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_800_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_800_inst_req_1 : boolean;
  signal type_cast_1054_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_800_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1084_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1301_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1075_inst_ack_1 : boolean;
  signal type_cast_804_inst_req_0 : boolean;
  signal type_cast_804_inst_ack_0 : boolean;
  signal type_cast_804_inst_req_1 : boolean;
  signal type_cast_804_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1066_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_818_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_818_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1081_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_818_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_818_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1289_inst_ack_0 : boolean;
  signal type_cast_822_inst_req_0 : boolean;
  signal type_cast_822_inst_ack_0 : boolean;
  signal type_cast_822_inst_req_1 : boolean;
  signal type_cast_822_inst_ack_1 : boolean;
  signal type_cast_1061_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1081_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1043_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1043_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1013_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1002_inst_ack_0 : boolean;
  signal ptr_deref_830_store_0_req_0 : boolean;
  signal WPIPE_Block0_start_1013_inst_req_1 : boolean;
  signal ptr_deref_830_store_0_ack_0 : boolean;
  signal WPIPE_Block1_start_1034_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_987_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1002_inst_req_0 : boolean;
  signal ptr_deref_830_store_0_req_1 : boolean;
  signal ptr_deref_830_store_0_ack_1 : boolean;
  signal type_cast_1338_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1013_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1013_inst_req_0 : boolean;
  signal WPIPE_Block0_start_987_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1034_inst_req_0 : boolean;
  signal if_stmt_844_branch_req_0 : boolean;
  signal if_stmt_844_branch_ack_1 : boolean;
  signal if_stmt_844_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_1072_inst_ack_1 : boolean;
  signal type_cast_855_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1043_inst_ack_0 : boolean;
  signal type_cast_855_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1072_inst_req_1 : boolean;
  signal type_cast_855_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1043_inst_req_0 : boolean;
  signal type_cast_855_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1078_inst_ack_1 : boolean;
  signal type_cast_1061_inst_req_1 : boolean;
  signal type_cast_859_inst_req_0 : boolean;
  signal type_cast_859_inst_ack_0 : boolean;
  signal type_cast_859_inst_req_1 : boolean;
  signal type_cast_859_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1078_inst_req_1 : boolean;
  signal type_cast_1061_inst_ack_0 : boolean;
  signal type_cast_863_inst_req_0 : boolean;
  signal type_cast_863_inst_ack_0 : boolean;
  signal type_cast_863_inst_req_1 : boolean;
  signal type_cast_863_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1066_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1072_inst_ack_0 : boolean;
  signal if_stmt_881_branch_req_0 : boolean;
  signal WPIPE_Block2_start_1075_inst_req_1 : boolean;
  signal if_stmt_881_branch_ack_1 : boolean;
  signal WPIPE_Block1_start_1031_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_984_inst_ack_1 : boolean;
  signal if_stmt_881_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_1031_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1081_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1289_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1072_inst_req_0 : boolean;
  signal type_cast_908_inst_req_0 : boolean;
  signal type_cast_908_inst_ack_0 : boolean;
  signal type_cast_908_inst_req_1 : boolean;
  signal type_cast_908_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1078_inst_ack_0 : boolean;
  signal type_cast_1426_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1081_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1069_inst_ack_0 : boolean;
  signal type_cast_1061_inst_req_0 : boolean;
  signal WPIPE_Block0_start_984_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1031_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1031_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1010_inst_ack_1 : boolean;
  signal array_obj_ref_937_index_offset_req_0 : boolean;
  signal WPIPE_Block1_start_1040_inst_ack_1 : boolean;
  signal array_obj_ref_937_index_offset_ack_0 : boolean;
  signal array_obj_ref_937_index_offset_req_1 : boolean;
  signal WPIPE_Block1_start_1040_inst_req_1 : boolean;
  signal array_obj_ref_937_index_offset_ack_1 : boolean;
  signal WPIPE_Block1_start_1069_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1010_inst_req_1 : boolean;
  signal addr_of_938_final_reg_req_0 : boolean;
  signal WPIPE_Block1_start_1040_inst_ack_0 : boolean;
  signal addr_of_938_final_reg_ack_0 : boolean;
  signal addr_of_938_final_reg_req_1 : boolean;
  signal WPIPE_Block1_start_1040_inst_req_0 : boolean;
  signal addr_of_938_final_reg_ack_1 : boolean;
  signal WPIPE_Block2_start_1078_inst_req_0 : boolean;
  signal ptr_deref_1372_load_0_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1301_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1010_inst_ack_0 : boolean;
  signal ptr_deref_941_store_0_req_0 : boolean;
  signal WPIPE_Block0_start_1010_inst_req_0 : boolean;
  signal ptr_deref_941_store_0_ack_0 : boolean;
  signal ptr_deref_941_store_0_req_1 : boolean;
  signal ptr_deref_941_store_0_ack_1 : boolean;
  signal WPIPE_Block2_start_1090_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1286_inst_req_1 : boolean;
  signal if_stmt_956_branch_req_0 : boolean;
  signal WPIPE_Block0_start_984_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_984_inst_req_0 : boolean;
  signal if_stmt_956_branch_ack_1 : boolean;
  signal if_stmt_956_branch_ack_0 : boolean;
  signal WPIPE_Block1_start_1028_inst_ack_1 : boolean;
  signal call_stmt_967_call_req_0 : boolean;
  signal call_stmt_967_call_ack_0 : boolean;
  signal type_cast_1446_inst_req_0 : boolean;
  signal call_stmt_967_call_req_1 : boolean;
  signal call_stmt_967_call_ack_1 : boolean;
  signal WPIPE_Block2_start_1087_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1093_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1298_inst_ack_1 : boolean;
  signal array_obj_ref_1367_index_offset_req_0 : boolean;
  signal WPIPE_Block1_start_1028_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1037_inst_ack_1 : boolean;
  signal type_cast_972_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1037_inst_req_1 : boolean;
  signal type_cast_972_inst_ack_0 : boolean;
  signal type_cast_972_inst_req_1 : boolean;
  signal type_cast_972_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_990_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1075_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1006_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_990_inst_req_1 : boolean;
  signal WPIPE_Block0_start_975_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1037_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_975_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_975_inst_req_1 : boolean;
  signal WPIPE_Block0_start_975_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1298_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1093_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1093_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1451_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1460_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1096_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1096_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1298_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1096_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1096_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1451_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1460_inst_req_0 : boolean;
  signal type_cast_1338_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1099_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1099_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1454_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1099_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1099_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1457_inst_ack_1 : boolean;
  signal type_cast_1386_inst_ack_1 : boolean;
  signal type_cast_1338_inst_req_0 : boolean;
  signal type_cast_1386_inst_req_1 : boolean;
  signal type_cast_1110_inst_req_0 : boolean;
  signal type_cast_1110_inst_ack_0 : boolean;
  signal type_cast_1110_inst_req_1 : boolean;
  signal ptr_deref_1372_load_0_ack_0 : boolean;
  signal type_cast_1110_inst_ack_1 : boolean;
  signal type_cast_1416_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1454_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1112_inst_req_0 : boolean;
  signal ptr_deref_1372_load_0_req_0 : boolean;
  signal WPIPE_Block2_start_1112_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1112_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1112_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1451_inst_ack_0 : boolean;
  signal type_cast_1386_inst_ack_0 : boolean;
  signal type_cast_1386_inst_req_0 : boolean;
  signal type_cast_1117_inst_req_0 : boolean;
  signal type_cast_1117_inst_ack_0 : boolean;
  signal type_cast_1117_inst_req_1 : boolean;
  signal type_cast_1117_inst_ack_1 : boolean;
  signal type_cast_1416_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1119_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1119_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1119_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1298_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1119_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1451_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1122_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1122_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1122_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1122_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1457_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1454_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1125_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1125_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1125_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1125_inst_ack_1 : boolean;
  signal type_cast_1416_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1454_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1128_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1128_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1128_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1128_inst_ack_1 : boolean;
  signal type_cast_1416_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1131_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1131_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1131_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1131_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1134_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1134_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1134_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1134_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1457_inst_ack_0 : boolean;
  signal type_cast_1376_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1137_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1137_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1137_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1137_inst_ack_1 : boolean;
  signal if_stmt_1311_branch_ack_0 : boolean;
  signal type_cast_1376_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1140_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1140_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1295_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1140_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1140_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1457_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1143_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1143_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1295_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1143_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1143_inst_ack_1 : boolean;
  signal if_stmt_1311_branch_ack_1 : boolean;
  signal WPIPE_Block3_start_1146_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1146_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1146_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1146_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1448_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1149_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1149_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1295_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1149_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1149_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1295_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1448_inst_req_1 : boolean;
  signal if_stmt_1311_branch_req_0 : boolean;
  signal type_cast_1406_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1152_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1152_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1152_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1152_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1448_inst_ack_0 : boolean;
  signal type_cast_1406_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1155_inst_req_0 : boolean;
  signal addr_of_1368_final_reg_ack_1 : boolean;
  signal WPIPE_Block3_start_1155_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1155_inst_req_1 : boolean;
  signal addr_of_1368_final_reg_req_1 : boolean;
  signal WPIPE_Block3_start_1155_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1448_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1307_inst_ack_1 : boolean;
  signal type_cast_1436_inst_ack_1 : boolean;
  signal type_cast_1166_inst_req_0 : boolean;
  signal type_cast_1166_inst_ack_0 : boolean;
  signal type_cast_1436_inst_req_1 : boolean;
  signal type_cast_1166_inst_req_1 : boolean;
  signal type_cast_1166_inst_ack_1 : boolean;
  signal type_cast_1376_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1307_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1168_inst_req_0 : boolean;
  signal addr_of_1368_final_reg_ack_0 : boolean;
  signal WPIPE_Block3_start_1168_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1292_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1168_inst_req_1 : boolean;
  signal addr_of_1368_final_reg_req_0 : boolean;
  signal WPIPE_Block3_start_1168_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1292_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1307_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1307_inst_req_0 : boolean;
  signal type_cast_1173_inst_req_0 : boolean;
  signal type_cast_1173_inst_ack_0 : boolean;
  signal type_cast_1173_inst_req_1 : boolean;
  signal type_cast_1173_inst_ack_1 : boolean;
  signal type_cast_1376_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1175_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1175_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1292_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1175_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1175_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1292_inst_req_0 : boolean;
  signal type_cast_1406_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1178_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1178_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1178_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1178_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1304_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1304_inst_req_1 : boolean;
  signal type_cast_1406_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1181_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1181_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1181_inst_req_1 : boolean;
  signal array_obj_ref_1367_index_offset_ack_1 : boolean;
  signal WPIPE_Block3_start_1181_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1184_inst_req_0 : boolean;
  signal array_obj_ref_1367_index_offset_req_1 : boolean;
  signal WPIPE_Block3_start_1184_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1184_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1184_inst_ack_1 : boolean;
  signal type_cast_1446_inst_ack_1 : boolean;
  signal type_cast_1446_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1304_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1304_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1188_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1188_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1289_inst_ack_1 : boolean;
  signal RPIPE_Block0_done_1188_inst_req_1 : boolean;
  signal array_obj_ref_1367_index_offset_ack_0 : boolean;
  signal RPIPE_Block0_done_1188_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1289_inst_req_1 : boolean;
  signal type_cast_1446_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1191_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1191_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1191_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1191_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1194_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1194_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1194_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1194_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1197_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1197_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1197_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1197_inst_ack_1 : boolean;
  signal call_stmt_1201_call_req_0 : boolean;
  signal call_stmt_1201_call_ack_0 : boolean;
  signal call_stmt_1201_call_req_1 : boolean;
  signal call_stmt_1201_call_ack_1 : boolean;
  signal type_cast_1205_inst_req_0 : boolean;
  signal type_cast_1205_inst_ack_0 : boolean;
  signal type_cast_1205_inst_req_1 : boolean;
  signal type_cast_1205_inst_ack_1 : boolean;
  signal type_cast_1214_inst_req_0 : boolean;
  signal type_cast_1214_inst_ack_0 : boolean;
  signal type_cast_1214_inst_req_1 : boolean;
  signal type_cast_1214_inst_ack_1 : boolean;
  signal type_cast_1224_inst_req_0 : boolean;
  signal type_cast_1224_inst_ack_0 : boolean;
  signal type_cast_1224_inst_req_1 : boolean;
  signal type_cast_1224_inst_ack_1 : boolean;
  signal type_cast_1234_inst_req_0 : boolean;
  signal type_cast_1234_inst_ack_0 : boolean;
  signal type_cast_1234_inst_req_1 : boolean;
  signal type_cast_1234_inst_ack_1 : boolean;
  signal type_cast_1436_inst_req_0 : boolean;
  signal type_cast_1244_inst_req_0 : boolean;
  signal type_cast_1244_inst_ack_0 : boolean;
  signal type_cast_1244_inst_req_1 : boolean;
  signal type_cast_1244_inst_ack_1 : boolean;
  signal type_cast_1254_inst_req_0 : boolean;
  signal type_cast_1254_inst_ack_0 : boolean;
  signal type_cast_1254_inst_req_1 : boolean;
  signal type_cast_1254_inst_ack_1 : boolean;
  signal type_cast_1264_inst_req_0 : boolean;
  signal type_cast_1264_inst_ack_0 : boolean;
  signal type_cast_1264_inst_req_1 : boolean;
  signal type_cast_1264_inst_ack_1 : boolean;
  signal type_cast_1274_inst_req_0 : boolean;
  signal type_cast_1274_inst_ack_0 : boolean;
  signal type_cast_1274_inst_req_1 : boolean;
  signal type_cast_1274_inst_ack_1 : boolean;
  signal type_cast_1284_inst_req_0 : boolean;
  signal type_cast_1284_inst_ack_0 : boolean;
  signal type_cast_1284_inst_req_1 : boolean;
  signal type_cast_1284_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1286_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1286_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1460_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1460_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1463_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1463_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1463_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1463_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1466_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1466_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1466_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1466_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1469_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1469_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1469_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1469_inst_ack_1 : boolean;
  signal if_stmt_1483_branch_req_0 : boolean;
  signal if_stmt_1483_branch_ack_1 : boolean;
  signal if_stmt_1483_branch_ack_0 : boolean;
  signal phi_stmt_474_req_0 : boolean;
  signal type_cast_480_inst_req_0 : boolean;
  signal type_cast_480_inst_ack_0 : boolean;
  signal type_cast_480_inst_req_1 : boolean;
  signal type_cast_480_inst_ack_1 : boolean;
  signal phi_stmt_474_req_1 : boolean;
  signal phi_stmt_474_ack_0 : boolean;
  signal phi_stmt_681_req_0 : boolean;
  signal type_cast_687_inst_req_0 : boolean;
  signal type_cast_687_inst_ack_0 : boolean;
  signal type_cast_687_inst_req_1 : boolean;
  signal type_cast_687_inst_ack_1 : boolean;
  signal phi_stmt_681_req_1 : boolean;
  signal phi_stmt_681_ack_0 : boolean;
  signal phi_stmt_925_req_1 : boolean;
  signal type_cast_928_inst_req_0 : boolean;
  signal type_cast_928_inst_ack_0 : boolean;
  signal type_cast_928_inst_req_1 : boolean;
  signal type_cast_928_inst_ack_1 : boolean;
  signal phi_stmt_925_req_0 : boolean;
  signal phi_stmt_925_ack_0 : boolean;
  signal phi_stmt_1355_req_0 : boolean;
  signal type_cast_1361_inst_req_0 : boolean;
  signal type_cast_1361_inst_ack_0 : boolean;
  signal type_cast_1361_inst_req_1 : boolean;
  signal type_cast_1361_inst_ack_1 : boolean;
  signal phi_stmt_1355_req_1 : boolean;
  signal phi_stmt_1355_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_34_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_34_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_34_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_34_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_34: Block -- control-path 
    signal convTranspose_CP_34_elements: BooleanArray(496 downto 0);
    -- 
  begin -- 
    convTranspose_CP_34_elements(0) <= convTranspose_CP_34_start;
    convTranspose_CP_34_symbol <= convTranspose_CP_34_elements(496);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	65 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	71 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	59 
    -- CP-element group 0: 	74 
    -- CP-element group 0: 	77 
    -- CP-element group 0: 	81 
    -- CP-element group 0: 	85 
    -- CP-element group 0: 	89 
    -- CP-element group 0: 	93 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	101 
    -- CP-element group 0: 	105 
    -- CP-element group 0: 	109 
    -- CP-element group 0: 	113 
    -- CP-element group 0: 	117 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0:  members (101) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_38/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/branch_block_stmt_38__entry__
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420__entry__
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_update_start_
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Update/cr
      -- 
    rr_130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => RPIPE_ConvTranspose_input_pipe_40_inst_req_0); -- 
    cr_149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_44_inst_req_1); -- 
    cr_177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_57_inst_req_1); -- 
    cr_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_69_inst_req_1); -- 
    cr_233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_82_inst_req_1); -- 
    cr_261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_94_inst_req_1); -- 
    cr_289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_107_inst_req_1); -- 
    cr_317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_119_inst_req_1); -- 
    cr_345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_132_inst_req_1); -- 
    cr_751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_345_inst_req_1); -- 
    cr_373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_144_inst_req_1); -- 
    cr_401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_157_inst_req_1); -- 
    cr_429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_169_inst_req_1); -- 
    cr_457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_182_inst_req_1); -- 
    cr_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_194_inst_req_1); -- 
    cr_513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_207_inst_req_1); -- 
    cr_527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_216_inst_req_1); -- 
    cr_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_220_inst_req_1); -- 
    cr_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_224_inst_req_1); -- 
    cr_569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_261_inst_req_1); -- 
    cr_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_265_inst_req_1); -- 
    cr_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_269_inst_req_1); -- 
    cr_611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_273_inst_req_1); -- 
    cr_639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_295_inst_req_1); -- 
    cr_667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_308_inst_req_1); -- 
    cr_695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_320_inst_req_1); -- 
    cr_723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_333_inst_req_1); -- 
    cr_779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_358_inst_req_1); -- 
    cr_807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_370_inst_req_1); -- 
    cr_835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_383_inst_req_1); -- 
    cr_863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_395_inst_req_1); -- 
    cr_891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(0), ack => type_cast_408_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_update_start_
      -- CP-element group 1: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Update/cr
      -- 
    ra_131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_40_inst_ack_0, ack => convTranspose_CP_34_elements(1)); -- 
    cr_135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(1), ack => RPIPE_ConvTranspose_input_pipe_40_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_40_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Sample/$entry
      -- 
    ca_136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_40_inst_ack_1, ack => convTranspose_CP_34_elements(2)); -- 
    rr_144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(2), ack => type_cast_44_inst_req_0); -- 
    rr_158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(2), ack => RPIPE_ConvTranspose_input_pipe_53_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Sample/ra
      -- 
    ra_145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_44_inst_ack_0, ack => convTranspose_CP_34_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	57 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_44_Update/ca
      -- 
    ca_150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_44_inst_ack_1, ack => convTranspose_CP_34_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_update_start_
      -- CP-element group 5: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Sample/$exit
      -- 
    ra_159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_53_inst_ack_0, ack => convTranspose_CP_34_elements(5)); -- 
    cr_163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(5), ack => RPIPE_ConvTranspose_input_pipe_53_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_53_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Sample/rr
      -- 
    ca_164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_53_inst_ack_1, ack => convTranspose_CP_34_elements(6)); -- 
    rr_172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(6), ack => type_cast_57_inst_req_0); -- 
    rr_186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(6), ack => RPIPE_ConvTranspose_input_pipe_65_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Sample/ra
      -- 
    ra_173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_57_inst_ack_0, ack => convTranspose_CP_34_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	57 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_57_Update/ca
      -- 
    ca_178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_57_inst_ack_1, ack => convTranspose_CP_34_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_update_start_
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Update/cr
      -- 
    ra_187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_65_inst_ack_0, ack => convTranspose_CP_34_elements(9)); -- 
    cr_191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(9), ack => RPIPE_ConvTranspose_input_pipe_65_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_65_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Sample/rr
      -- 
    ca_192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_65_inst_ack_1, ack => convTranspose_CP_34_elements(10)); -- 
    rr_200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(10), ack => type_cast_69_inst_req_0); -- 
    rr_214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(10), ack => RPIPE_ConvTranspose_input_pipe_78_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Sample/ra
      -- 
    ra_201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_69_inst_ack_0, ack => convTranspose_CP_34_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	60 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_69_Update/ca
      -- 
    ca_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_69_inst_ack_1, ack => convTranspose_CP_34_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_update_start_
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Update/cr
      -- 
    ra_215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_78_inst_ack_0, ack => convTranspose_CP_34_elements(13)); -- 
    cr_219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(13), ack => RPIPE_ConvTranspose_input_pipe_78_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_78_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Sample/rr
      -- 
    ca_220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_78_inst_ack_1, ack => convTranspose_CP_34_elements(14)); -- 
    rr_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(14), ack => type_cast_82_inst_req_0); -- 
    rr_242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(14), ack => RPIPE_ConvTranspose_input_pipe_90_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Sample/ra
      -- 
    ra_229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_82_inst_ack_0, ack => convTranspose_CP_34_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	60 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_82_Update/ca
      -- 
    ca_234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_82_inst_ack_1, ack => convTranspose_CP_34_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_update_start_
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Update/cr
      -- 
    ra_243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_90_inst_ack_0, ack => convTranspose_CP_34_elements(17)); -- 
    cr_247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(17), ack => RPIPE_ConvTranspose_input_pipe_90_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_90_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Sample/rr
      -- 
    ca_248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_90_inst_ack_1, ack => convTranspose_CP_34_elements(18)); -- 
    rr_256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(18), ack => type_cast_94_inst_req_0); -- 
    rr_270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(18), ack => RPIPE_ConvTranspose_input_pipe_103_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Sample/ra
      -- 
    ra_257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_94_inst_ack_0, ack => convTranspose_CP_34_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	63 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_94_Update/ca
      -- 
    ca_262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_94_inst_ack_1, ack => convTranspose_CP_34_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_update_start_
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Update/cr
      -- 
    ra_271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_103_inst_ack_0, ack => convTranspose_CP_34_elements(21)); -- 
    cr_275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(21), ack => RPIPE_ConvTranspose_input_pipe_103_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_103_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Sample/rr
      -- 
    ca_276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_103_inst_ack_1, ack => convTranspose_CP_34_elements(22)); -- 
    rr_284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(22), ack => type_cast_107_inst_req_0); -- 
    rr_298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(22), ack => RPIPE_ConvTranspose_input_pipe_115_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Sample/ra
      -- 
    ra_285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_107_inst_ack_0, ack => convTranspose_CP_34_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	63 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_107_Update/ca
      -- 
    ca_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_107_inst_ack_1, ack => convTranspose_CP_34_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_update_start_
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Update/cr
      -- 
    ra_299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_115_inst_ack_0, ack => convTranspose_CP_34_elements(25)); -- 
    cr_303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(25), ack => RPIPE_ConvTranspose_input_pipe_115_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_115_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Sample/rr
      -- 
    ca_304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_115_inst_ack_1, ack => convTranspose_CP_34_elements(26)); -- 
    rr_312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(26), ack => type_cast_119_inst_req_0); -- 
    rr_326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(26), ack => RPIPE_ConvTranspose_input_pipe_128_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Sample/ra
      -- 
    ra_313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_119_inst_ack_0, ack => convTranspose_CP_34_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	66 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_119_Update/ca
      -- 
    ca_318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_119_inst_ack_1, ack => convTranspose_CP_34_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_update_start_
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Update/cr
      -- 
    ra_327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_128_inst_ack_0, ack => convTranspose_CP_34_elements(29)); -- 
    cr_331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(29), ack => RPIPE_ConvTranspose_input_pipe_128_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_128_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Sample/rr
      -- 
    ca_332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_128_inst_ack_1, ack => convTranspose_CP_34_elements(30)); -- 
    rr_340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(30), ack => type_cast_132_inst_req_0); -- 
    rr_354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(30), ack => RPIPE_ConvTranspose_input_pipe_140_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Sample/ra
      -- 
    ra_341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_132_inst_ack_0, ack => convTranspose_CP_34_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	66 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_132_Update/ca
      -- 
    ca_346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_132_inst_ack_1, ack => convTranspose_CP_34_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_update_start_
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Update/cr
      -- 
    ra_355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_140_inst_ack_0, ack => convTranspose_CP_34_elements(33)); -- 
    cr_359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(33), ack => RPIPE_ConvTranspose_input_pipe_140_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_140_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Sample/rr
      -- 
    ca_360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_140_inst_ack_1, ack => convTranspose_CP_34_elements(34)); -- 
    rr_368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(34), ack => type_cast_144_inst_req_0); -- 
    rr_382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(34), ack => RPIPE_ConvTranspose_input_pipe_153_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Sample/ra
      -- 
    ra_369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_144_inst_ack_0, ack => convTranspose_CP_34_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	69 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_144_Update/ca
      -- 
    ca_374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_144_inst_ack_1, ack => convTranspose_CP_34_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_update_start_
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Update/cr
      -- 
    ra_383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_153_inst_ack_0, ack => convTranspose_CP_34_elements(37)); -- 
    cr_387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(37), ack => RPIPE_ConvTranspose_input_pipe_153_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_153_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Sample/rr
      -- 
    ca_388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_153_inst_ack_1, ack => convTranspose_CP_34_elements(38)); -- 
    rr_396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(38), ack => type_cast_157_inst_req_0); -- 
    rr_410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(38), ack => RPIPE_ConvTranspose_input_pipe_165_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Sample/ra
      -- 
    ra_397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_157_inst_ack_0, ack => convTranspose_CP_34_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	69 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_157_Update/ca
      -- 
    ca_402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_157_inst_ack_1, ack => convTranspose_CP_34_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_update_start_
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Update/cr
      -- 
    ra_411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_165_inst_ack_0, ack => convTranspose_CP_34_elements(41)); -- 
    cr_415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(41), ack => RPIPE_ConvTranspose_input_pipe_165_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_165_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Sample/rr
      -- 
    ca_416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_165_inst_ack_1, ack => convTranspose_CP_34_elements(42)); -- 
    rr_424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(42), ack => type_cast_169_inst_req_0); -- 
    rr_438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(42), ack => RPIPE_ConvTranspose_input_pipe_178_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Sample/ra
      -- 
    ra_425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_169_inst_ack_0, ack => convTranspose_CP_34_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	72 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_169_Update/ca
      -- 
    ca_430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_169_inst_ack_1, ack => convTranspose_CP_34_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_update_start_
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Update/cr
      -- 
    ra_439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_178_inst_ack_0, ack => convTranspose_CP_34_elements(45)); -- 
    cr_443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(45), ack => RPIPE_ConvTranspose_input_pipe_178_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_178_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Sample/rr
      -- 
    ca_444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_178_inst_ack_1, ack => convTranspose_CP_34_elements(46)); -- 
    rr_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(46), ack => RPIPE_ConvTranspose_input_pipe_190_inst_req_0); -- 
    rr_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(46), ack => type_cast_182_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Sample/ra
      -- 
    ra_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_182_inst_ack_0, ack => convTranspose_CP_34_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	72 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_182_Update/ca
      -- 
    ca_458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_182_inst_ack_1, ack => convTranspose_CP_34_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_update_start_
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Update/cr
      -- 
    ra_467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_190_inst_ack_0, ack => convTranspose_CP_34_elements(49)); -- 
    cr_471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(49), ack => RPIPE_ConvTranspose_input_pipe_190_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_190_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Sample/rr
      -- 
    ca_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_190_inst_ack_1, ack => convTranspose_CP_34_elements(50)); -- 
    rr_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(50), ack => type_cast_194_inst_req_0); -- 
    rr_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(50), ack => RPIPE_ConvTranspose_input_pipe_203_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Sample/ra
      -- 
    ra_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_194_inst_ack_0, ack => convTranspose_CP_34_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	75 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_194_Update/ca
      -- 
    ca_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_194_inst_ack_1, ack => convTranspose_CP_34_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_update_start_
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Update/cr
      -- 
    ra_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_203_inst_ack_0, ack => convTranspose_CP_34_elements(53)); -- 
    cr_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(53), ack => RPIPE_ConvTranspose_input_pipe_203_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	78 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_203_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Sample/rr
      -- 
    ca_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_203_inst_ack_1, ack => convTranspose_CP_34_elements(54)); -- 
    rr_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(54), ack => type_cast_207_inst_req_0); -- 
    rr_620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(54), ack => RPIPE_ConvTranspose_input_pipe_291_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Sample/ra
      -- 
    ra_509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_207_inst_ack_0, ack => convTranspose_CP_34_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	75 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_207_Update/ca
      -- 
    ca_514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_207_inst_ack_1, ack => convTranspose_CP_34_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	4 
    -- CP-element group 57: 	8 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Sample/rr
      -- 
    rr_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(57), ack => type_cast_216_inst_req_0); -- 
    convTranspose_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(4) & convTranspose_CP_34_elements(8);
      gj_convTranspose_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Sample/ra
      -- 
    ra_523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_216_inst_ack_0, ack => convTranspose_CP_34_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	0 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	118 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_216_Update/ca
      -- 
    ca_528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_216_inst_ack_1, ack => convTranspose_CP_34_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	12 
    -- CP-element group 60: 	16 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Sample/rr
      -- 
    rr_536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(60), ack => type_cast_220_inst_req_0); -- 
    convTranspose_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(12) & convTranspose_CP_34_elements(16);
      gj_convTranspose_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Sample/ra
      -- 
    ra_537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_220_inst_ack_0, ack => convTranspose_CP_34_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	118 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_220_Update/ca
      -- 
    ca_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_220_inst_ack_1, ack => convTranspose_CP_34_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	20 
    -- CP-element group 63: 	24 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Sample/rr
      -- 
    rr_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(63), ack => type_cast_224_inst_req_0); -- 
    convTranspose_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(20) & convTranspose_CP_34_elements(24);
      gj_convTranspose_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Sample/ra
      -- 
    ra_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_224_inst_ack_0, ack => convTranspose_CP_34_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	0 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	118 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_224_Update/ca
      -- 
    ca_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_224_inst_ack_1, ack => convTranspose_CP_34_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	28 
    -- CP-element group 66: 	32 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Sample/rr
      -- 
    rr_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(66), ack => type_cast_261_inst_req_0); -- 
    convTranspose_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(28) & convTranspose_CP_34_elements(32);
      gj_convTranspose_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Sample/ra
      -- 
    ra_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_261_inst_ack_0, ack => convTranspose_CP_34_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	118 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_261_Update/ca
      -- 
    ca_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_261_inst_ack_1, ack => convTranspose_CP_34_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	40 
    -- CP-element group 69: 	36 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Sample/rr
      -- 
    rr_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(69), ack => type_cast_265_inst_req_0); -- 
    convTranspose_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(40) & convTranspose_CP_34_elements(36);
      gj_convTranspose_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Sample/ra
      -- 
    ra_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_265_inst_ack_0, ack => convTranspose_CP_34_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	0 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	118 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_265_Update/ca
      -- 
    ca_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_265_inst_ack_1, ack => convTranspose_CP_34_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	44 
    -- CP-element group 72: 	48 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Sample/rr
      -- 
    rr_592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(72), ack => type_cast_269_inst_req_0); -- 
    convTranspose_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(44) & convTranspose_CP_34_elements(48);
      gj_convTranspose_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Sample/ra
      -- 
    ra_593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_269_inst_ack_0, ack => convTranspose_CP_34_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	0 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	118 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_269_Update/ca
      -- 
    ca_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_269_inst_ack_1, ack => convTranspose_CP_34_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	56 
    -- CP-element group 75: 	52 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Sample/rr
      -- 
    rr_606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(75), ack => type_cast_273_inst_req_0); -- 
    convTranspose_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(56) & convTranspose_CP_34_elements(52);
      gj_convTranspose_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Sample/ra
      -- 
    ra_607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_273_inst_ack_0, ack => convTranspose_CP_34_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	0 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	118 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_273_Update/ca
      -- 
    ca_612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_273_inst_ack_1, ack => convTranspose_CP_34_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	54 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_update_start_
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Update/cr
      -- 
    ra_621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_291_inst_ack_0, ack => convTranspose_CP_34_elements(78)); -- 
    cr_625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(78), ack => RPIPE_ConvTranspose_input_pipe_291_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_291_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Sample/rr
      -- 
    ca_626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_291_inst_ack_1, ack => convTranspose_CP_34_elements(79)); -- 
    rr_634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(79), ack => type_cast_295_inst_req_0); -- 
    rr_648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(79), ack => RPIPE_ConvTranspose_input_pipe_304_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Sample/ra
      -- 
    ra_635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_295_inst_ack_0, ack => convTranspose_CP_34_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	0 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	118 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_295_Update/ca
      -- 
    ca_640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_295_inst_ack_1, ack => convTranspose_CP_34_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_update_start_
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Update/cr
      -- 
    ra_649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_304_inst_ack_0, ack => convTranspose_CP_34_elements(82)); -- 
    cr_653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(82), ack => RPIPE_ConvTranspose_input_pipe_304_inst_req_1); -- 
    -- CP-element group 83:  fork  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_304_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Sample/rr
      -- 
    ca_654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_304_inst_ack_1, ack => convTranspose_CP_34_elements(83)); -- 
    rr_662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(83), ack => type_cast_308_inst_req_0); -- 
    rr_676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(83), ack => RPIPE_ConvTranspose_input_pipe_316_inst_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Sample/ra
      -- 
    ra_663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_308_inst_ack_0, ack => convTranspose_CP_34_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	0 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	118 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_308_Update/ca
      -- 
    ca_668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_308_inst_ack_1, ack => convTranspose_CP_34_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_update_start_
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Update/cr
      -- 
    ra_677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_316_inst_ack_0, ack => convTranspose_CP_34_elements(86)); -- 
    cr_681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(86), ack => RPIPE_ConvTranspose_input_pipe_316_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_316_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Sample/rr
      -- 
    ca_682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_316_inst_ack_1, ack => convTranspose_CP_34_elements(87)); -- 
    rr_690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(87), ack => type_cast_320_inst_req_0); -- 
    rr_704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(87), ack => RPIPE_ConvTranspose_input_pipe_329_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Sample/ra
      -- 
    ra_691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_320_inst_ack_0, ack => convTranspose_CP_34_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	0 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	118 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_320_Update/ca
      -- 
    ca_696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_320_inst_ack_1, ack => convTranspose_CP_34_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_update_start_
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Update/cr
      -- 
    ra_705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_329_inst_ack_0, ack => convTranspose_CP_34_elements(90)); -- 
    cr_709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(90), ack => RPIPE_ConvTranspose_input_pipe_329_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_329_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Sample/rr
      -- 
    ca_710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_329_inst_ack_1, ack => convTranspose_CP_34_elements(91)); -- 
    rr_718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(91), ack => type_cast_333_inst_req_0); -- 
    rr_732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(91), ack => RPIPE_ConvTranspose_input_pipe_341_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Sample/ra
      -- 
    ra_719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_333_inst_ack_0, ack => convTranspose_CP_34_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	0 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	118 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_333_Update/ca
      -- 
    ca_724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_333_inst_ack_1, ack => convTranspose_CP_34_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_update_start_
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Update/cr
      -- 
    ra_733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_341_inst_ack_0, ack => convTranspose_CP_34_elements(94)); -- 
    cr_737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(94), ack => RPIPE_ConvTranspose_input_pipe_341_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_341_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Sample/rr
      -- 
    ca_738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_341_inst_ack_1, ack => convTranspose_CP_34_elements(95)); -- 
    rr_746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(95), ack => type_cast_345_inst_req_0); -- 
    rr_760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(95), ack => RPIPE_ConvTranspose_input_pipe_354_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Sample/ra
      -- 
    ra_747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_345_inst_ack_0, ack => convTranspose_CP_34_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	118 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_345_Update/$exit
      -- 
    ca_752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_345_inst_ack_1, ack => convTranspose_CP_34_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_update_start_
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Update/cr
      -- 
    ra_761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_354_inst_ack_0, ack => convTranspose_CP_34_elements(98)); -- 
    cr_765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(98), ack => RPIPE_ConvTranspose_input_pipe_354_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_354_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Sample/rr
      -- 
    ca_766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_354_inst_ack_1, ack => convTranspose_CP_34_elements(99)); -- 
    rr_774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(99), ack => type_cast_358_inst_req_0); -- 
    rr_788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(99), ack => RPIPE_ConvTranspose_input_pipe_366_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Sample/ra
      -- 
    ra_775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_358_inst_ack_0, ack => convTranspose_CP_34_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	0 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	118 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_358_Update/ca
      -- 
    ca_780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_358_inst_ack_1, ack => convTranspose_CP_34_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_update_start_
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Update/cr
      -- 
    ra_789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_366_inst_ack_0, ack => convTranspose_CP_34_elements(102)); -- 
    cr_793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(102), ack => RPIPE_ConvTranspose_input_pipe_366_inst_req_1); -- 
    -- CP-element group 103:  fork  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_366_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Sample/rr
      -- 
    ca_794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_366_inst_ack_1, ack => convTranspose_CP_34_elements(103)); -- 
    rr_802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(103), ack => type_cast_370_inst_req_0); -- 
    rr_816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(103), ack => RPIPE_ConvTranspose_input_pipe_379_inst_req_0); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Sample/ra
      -- 
    ra_803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_370_inst_ack_0, ack => convTranspose_CP_34_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	0 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	118 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_370_Update/ca
      -- 
    ca_808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_370_inst_ack_1, ack => convTranspose_CP_34_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_update_start_
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Update/cr
      -- 
    ra_817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_379_inst_ack_0, ack => convTranspose_CP_34_elements(106)); -- 
    cr_821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(106), ack => RPIPE_ConvTranspose_input_pipe_379_inst_req_1); -- 
    -- CP-element group 107:  fork  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_379_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Sample/rr
      -- 
    ca_822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_379_inst_ack_1, ack => convTranspose_CP_34_elements(107)); -- 
    rr_830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(107), ack => type_cast_383_inst_req_0); -- 
    rr_844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(107), ack => RPIPE_ConvTranspose_input_pipe_391_inst_req_0); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Sample/ra
      -- 
    ra_831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_383_inst_ack_0, ack => convTranspose_CP_34_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	0 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	118 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_383_Update/ca
      -- 
    ca_836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_383_inst_ack_1, ack => convTranspose_CP_34_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_update_start_
      -- CP-element group 110: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Update/cr
      -- 
    ra_845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_391_inst_ack_0, ack => convTranspose_CP_34_elements(110)); -- 
    cr_849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(110), ack => RPIPE_ConvTranspose_input_pipe_391_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_391_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Sample/rr
      -- 
    ca_850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_391_inst_ack_1, ack => convTranspose_CP_34_elements(111)); -- 
    rr_858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(111), ack => type_cast_395_inst_req_0); -- 
    rr_872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(111), ack => RPIPE_ConvTranspose_input_pipe_404_inst_req_0); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Sample/ra
      -- 
    ra_859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_395_inst_ack_0, ack => convTranspose_CP_34_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	0 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	118 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_395_Update/ca
      -- 
    ca_864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_395_inst_ack_1, ack => convTranspose_CP_34_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_update_start_
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Update/cr
      -- 
    ra_873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_404_inst_ack_0, ack => convTranspose_CP_34_elements(114)); -- 
    cr_877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(114), ack => RPIPE_ConvTranspose_input_pipe_404_inst_req_1); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/RPIPE_ConvTranspose_input_pipe_404_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Sample/rr
      -- 
    ca_878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_404_inst_ack_1, ack => convTranspose_CP_34_elements(115)); -- 
    rr_886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(115), ack => type_cast_408_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Sample/ra
      -- 
    ra_887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_408_inst_ack_0, ack => convTranspose_CP_34_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	0 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/type_cast_408_Update/ca
      -- 
    ca_892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_408_inst_ack_1, ack => convTranspose_CP_34_elements(117)); -- 
    -- CP-element group 118:  branch  join  transition  place  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	62 
    -- CP-element group 118: 	65 
    -- CP-element group 118: 	68 
    -- CP-element group 118: 	71 
    -- CP-element group 118: 	59 
    -- CP-element group 118: 	74 
    -- CP-element group 118: 	77 
    -- CP-element group 118: 	81 
    -- CP-element group 118: 	85 
    -- CP-element group 118: 	89 
    -- CP-element group 118: 	93 
    -- CP-element group 118: 	97 
    -- CP-element group 118: 	101 
    -- CP-element group 118: 	105 
    -- CP-element group 118: 	109 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (10) 
      -- CP-element group 118: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420__exit__
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421__entry__
      -- CP-element group 118: 	 branch_block_stmt_38/assign_stmt_41_to_assign_stmt_420/$exit
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421_dead_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421_eval_test/$entry
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421_eval_test/$exit
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421_eval_test/branch_req
      -- CP-element group 118: 	 branch_block_stmt_38/R_cmp513_422_place
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421_if_link/$entry
      -- CP-element group 118: 	 branch_block_stmt_38/if_stmt_421_else_link/$entry
      -- 
    branch_req_900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(118), ack => if_stmt_421_branch_req_0); -- 
    convTranspose_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(62) & convTranspose_CP_34_elements(65) & convTranspose_CP_34_elements(68) & convTranspose_CP_34_elements(71) & convTranspose_CP_34_elements(59) & convTranspose_CP_34_elements(74) & convTranspose_CP_34_elements(77) & convTranspose_CP_34_elements(81) & convTranspose_CP_34_elements(85) & convTranspose_CP_34_elements(89) & convTranspose_CP_34_elements(93) & convTranspose_CP_34_elements(97) & convTranspose_CP_34_elements(101) & convTranspose_CP_34_elements(105) & convTranspose_CP_34_elements(109) & convTranspose_CP_34_elements(113) & convTranspose_CP_34_elements(117);
      gj_convTranspose_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	123 
    -- CP-element group 119: 	124 
    -- CP-element group 119:  members (18) 
      -- CP-element group 119: 	 branch_block_stmt_38/merge_stmt_442__exit__
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471__entry__
      -- CP-element group 119: 	 branch_block_stmt_38/if_stmt_421_if_link/$exit
      -- CP-element group 119: 	 branch_block_stmt_38/if_stmt_421_if_link/if_choice_transition
      -- CP-element group 119: 	 branch_block_stmt_38/entry_bbx_xnph515
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_update_start_
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_38/entry_bbx_xnph515_PhiReq/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/entry_bbx_xnph515_PhiReq/$exit
      -- CP-element group 119: 	 branch_block_stmt_38/merge_stmt_442_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_38/merge_stmt_442_PhiAck/$entry
      -- CP-element group 119: 	 branch_block_stmt_38/merge_stmt_442_PhiAck/$exit
      -- CP-element group 119: 	 branch_block_stmt_38/merge_stmt_442_PhiAck/dummy
      -- 
    if_choice_transition_905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_421_branch_ack_1, ack => convTranspose_CP_34_elements(119)); -- 
    rr_944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(119), ack => type_cast_457_inst_req_0); -- 
    cr_949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(119), ack => type_cast_457_inst_req_1); -- 
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	469 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_38/if_stmt_421_else_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_38/if_stmt_421_else_link/else_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_38/entry_forx_xcond190x_xpreheader
      -- CP-element group 120: 	 branch_block_stmt_38/entry_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 120: 	 branch_block_stmt_38/entry_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_421_branch_ack_0, ack => convTranspose_CP_34_elements(120)); -- 
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	469 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	167 
    -- CP-element group 121: 	168 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_38/merge_stmt_643__exit__
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678__entry__
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_update_start_
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/if_stmt_436_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_38/if_stmt_436_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xcond190x_xpreheader_bbx_xnph511
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xcond190x_xpreheader_bbx_xnph511_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/forx_xcond190x_xpreheader_bbx_xnph511_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_38/merge_stmt_643_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_38/merge_stmt_643_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_38/merge_stmt_643_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_38/merge_stmt_643_PhiAck/dummy
      -- 
    if_choice_transition_927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_436_branch_ack_1, ack => convTranspose_CP_34_elements(121)); -- 
    cr_1308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(121), ack => type_cast_664_inst_req_1); -- 
    rr_1303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(121), ack => type_cast_664_inst_req_0); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	469 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	482 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_38/if_stmt_436_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_38/if_stmt_436_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_38/forx_xcond190x_xpreheader_forx_xend250
      -- CP-element group 122: 	 branch_block_stmt_38/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_38/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$exit
      -- 
    else_choice_transition_931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_436_branch_ack_0, ack => convTranspose_CP_34_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	119 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Sample/ra
      -- 
    ra_945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_457_inst_ack_0, ack => convTranspose_CP_34_elements(123)); -- 
    -- CP-element group 124:  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	119 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	470 
    -- CP-element group 124:  members (9) 
      -- CP-element group 124: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471__exit__
      -- CP-element group 124: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody
      -- CP-element group 124: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/$exit
      -- CP-element group 124: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_38/assign_stmt_448_to_assign_stmt_471/type_cast_457_Update/ca
      -- CP-element group 124: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/$entry
      -- CP-element group 124: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_474/$entry
      -- CP-element group 124: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/$entry
      -- 
    ca_950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_457_inst_ack_1, ack => convTranspose_CP_34_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	475 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	164 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_sample_complete
      -- CP-element group 125: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Sample/ack
      -- 
    ack_979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_486_index_offset_ack_0, ack => convTranspose_CP_34_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	475 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (11) 
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_root_address_calculated
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_offset_calculated
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Update/ack
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_base_plus_offset/$entry
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_base_plus_offset/$exit
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_base_plus_offset/sum_rename_req
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_base_plus_offset/sum_rename_ack
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_request/$entry
      -- CP-element group 126: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_request/req
      -- 
    ack_984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_486_index_offset_ack_1, ack => convTranspose_CP_34_elements(126)); -- 
    req_993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(126), ack => addr_of_487_final_reg_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_request/$exit
      -- CP-element group 127: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_request/ack
      -- 
    ack_994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_487_final_reg_ack_0, ack => convTranspose_CP_34_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	475 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	161 
    -- CP-element group 128:  members (19) 
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_word_addrgen/root_register_ack
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_word_addrgen/root_register_req
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_word_addrgen/$exit
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_word_addrgen/$entry
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_plus_offset/sum_rename_ack
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_plus_offset/sum_rename_req
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_plus_offset/$exit
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_plus_offset/$entry
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_addr_resize/base_resize_ack
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_addr_resize/base_resize_req
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_addr_resize/$exit
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_addr_resize/$entry
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_address_resized
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_root_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_word_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_base_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_complete/$exit
      -- CP-element group 128: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_complete/ack
      -- 
    ack_999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_487_final_reg_ack_1, ack => convTranspose_CP_34_elements(128)); -- 
    -- CP-element group 129:  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	475 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (6) 
      -- CP-element group 129: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_update_start_
      -- CP-element group 129: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Update/$entry
      -- CP-element group 129: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Update/cr
      -- 
    ra_1008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_490_inst_ack_0, ack => convTranspose_CP_34_elements(129)); -- 
    cr_1012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(129), ack => RPIPE_ConvTranspose_input_pipe_490_inst_req_1); -- 
    -- CP-element group 130:  fork  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: 	133 
    -- CP-element group 130:  members (9) 
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Sample/rr
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Sample/rr
      -- 
    ca_1013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_490_inst_ack_1, ack => convTranspose_CP_34_elements(130)); -- 
    rr_1021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(130), ack => type_cast_494_inst_req_0); -- 
    rr_1035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(130), ack => RPIPE_ConvTranspose_input_pipe_503_inst_req_0); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Sample/ra
      -- 
    ra_1022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_494_inst_ack_0, ack => convTranspose_CP_34_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	475 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	161 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Update/ca
      -- 
    ca_1027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_494_inst_ack_1, ack => convTranspose_CP_34_elements(132)); -- 
    -- CP-element group 133:  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	130 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_update_start_
      -- CP-element group 133: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Update/cr
      -- 
    ra_1036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_503_inst_ack_0, ack => convTranspose_CP_34_elements(133)); -- 
    cr_1040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(133), ack => RPIPE_ConvTranspose_input_pipe_503_inst_req_1); -- 
    -- CP-element group 134:  fork  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (9) 
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_503_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Sample/rr
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Sample/rr
      -- 
    ca_1041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_503_inst_ack_1, ack => convTranspose_CP_34_elements(134)); -- 
    rr_1049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(134), ack => type_cast_507_inst_req_0); -- 
    rr_1063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(134), ack => RPIPE_ConvTranspose_input_pipe_521_inst_req_0); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Sample/ra
      -- 
    ra_1050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_507_inst_ack_0, ack => convTranspose_CP_34_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	475 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	161 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Update/ca
      -- 
    ca_1055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_507_inst_ack_1, ack => convTranspose_CP_34_elements(136)); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_update_start_
      -- CP-element group 137: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Update/cr
      -- 
    ra_1064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_521_inst_ack_0, ack => convTranspose_CP_34_elements(137)); -- 
    cr_1068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(137), ack => RPIPE_ConvTranspose_input_pipe_521_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138: 	141 
    -- CP-element group 138:  members (9) 
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_521_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_sample_start_
      -- 
    ca_1069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_521_inst_ack_1, ack => convTranspose_CP_34_elements(138)); -- 
    rr_1077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(138), ack => type_cast_525_inst_req_0); -- 
    rr_1091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(138), ack => RPIPE_ConvTranspose_input_pipe_539_inst_req_0); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Sample/ra
      -- 
    ra_1078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_525_inst_ack_0, ack => convTranspose_CP_34_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	475 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	161 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Update/ca
      -- 
    ca_1083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_525_inst_ack_1, ack => convTranspose_CP_34_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	138 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (6) 
      -- CP-element group 141: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Update/cr
      -- CP-element group 141: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Update/$entry
      -- CP-element group 141: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_update_start_
      -- 
    ra_1092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_539_inst_ack_0, ack => convTranspose_CP_34_elements(141)); -- 
    cr_1096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(141), ack => RPIPE_ConvTranspose_input_pipe_539_inst_req_1); -- 
    -- CP-element group 142:  fork  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	145 
    -- CP-element group 142:  members (9) 
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_539_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Sample/rr
      -- CP-element group 142: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Sample/$entry
      -- 
    ca_1097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_539_inst_ack_1, ack => convTranspose_CP_34_elements(142)); -- 
    rr_1105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(142), ack => type_cast_543_inst_req_0); -- 
    rr_1119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(142), ack => RPIPE_ConvTranspose_input_pipe_557_inst_req_0); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Sample/$exit
      -- 
    ra_1106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_543_inst_ack_0, ack => convTranspose_CP_34_elements(143)); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	475 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	161 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Update/$exit
      -- 
    ca_1111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_543_inst_ack_1, ack => convTranspose_CP_34_elements(144)); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	142 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_update_start_
      -- CP-element group 145: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Sample/ra
      -- 
    ra_1120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_557_inst_ack_0, ack => convTranspose_CP_34_elements(145)); -- 
    cr_1124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(145), ack => RPIPE_ConvTranspose_input_pipe_557_inst_req_1); -- 
    -- CP-element group 146:  fork  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	149 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Sample/rr
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Update/ca
      -- CP-element group 146: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_557_Update/$exit
      -- 
    ca_1125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_557_inst_ack_1, ack => convTranspose_CP_34_elements(146)); -- 
    rr_1133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(146), ack => type_cast_561_inst_req_0); -- 
    rr_1147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(146), ack => RPIPE_ConvTranspose_input_pipe_575_inst_req_0); -- 
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_sample_completed_
      -- 
    ra_1134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_561_inst_ack_0, ack => convTranspose_CP_34_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	475 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	161 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_update_completed_
      -- 
    ca_1139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_561_inst_ack_1, ack => convTranspose_CP_34_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	146 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (6) 
      -- CP-element group 149: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Update/$entry
      -- CP-element group 149: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Sample/ra
      -- CP-element group 149: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_update_start_
      -- CP-element group 149: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_sample_completed_
      -- 
    ra_1148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_575_inst_ack_0, ack => convTranspose_CP_34_elements(149)); -- 
    cr_1152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(149), ack => RPIPE_ConvTranspose_input_pipe_575_inst_req_1); -- 
    -- CP-element group 150:  fork  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (9) 
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Update/ca
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_575_update_completed_
      -- 
    ca_1153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_575_inst_ack_1, ack => convTranspose_CP_34_elements(150)); -- 
    rr_1161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(150), ack => type_cast_579_inst_req_0); -- 
    rr_1175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(150), ack => RPIPE_ConvTranspose_input_pipe_593_inst_req_0); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_sample_completed_
      -- 
    ra_1162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_579_inst_ack_0, ack => convTranspose_CP_34_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	475 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	161 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_update_completed_
      -- 
    ca_1167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_579_inst_ack_1, ack => convTranspose_CP_34_elements(152)); -- 
    -- CP-element group 153:  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	150 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (6) 
      -- CP-element group 153: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Sample/ra
      -- CP-element group 153: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_update_start_
      -- CP-element group 153: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_sample_completed_
      -- 
    ra_1176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_593_inst_ack_0, ack => convTranspose_CP_34_elements(153)); -- 
    cr_1180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(153), ack => RPIPE_ConvTranspose_input_pipe_593_inst_req_1); -- 
    -- CP-element group 154:  fork  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	157 
    -- CP-element group 154:  members (9) 
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Update/ca
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_593_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_sample_start_
      -- 
    ca_1181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_593_inst_ack_1, ack => convTranspose_CP_34_elements(154)); -- 
    rr_1189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(154), ack => type_cast_597_inst_req_0); -- 
    rr_1203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(154), ack => RPIPE_ConvTranspose_input_pipe_611_inst_req_0); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Sample/$exit
      -- 
    ra_1190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_597_inst_ack_0, ack => convTranspose_CP_34_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	475 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	161 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Update/ca
      -- CP-element group 156: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_update_completed_
      -- 
    ca_1195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_597_inst_ack_1, ack => convTranspose_CP_34_elements(156)); -- 
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Update/cr
      -- CP-element group 157: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Sample/ra
      -- CP-element group 157: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_update_start_
      -- CP-element group 157: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_sample_completed_
      -- 
    ra_1204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_611_inst_ack_0, ack => convTranspose_CP_34_elements(157)); -- 
    cr_1208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(157), ack => RPIPE_ConvTranspose_input_pipe_611_inst_req_1); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Sample/rr
      -- CP-element group 158: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Update/ca
      -- CP-element group 158: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_611_update_completed_
      -- 
    ca_1209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_611_inst_ack_1, ack => convTranspose_CP_34_elements(158)); -- 
    rr_1217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(158), ack => type_cast_615_inst_req_0); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Sample/ra
      -- CP-element group 159: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_sample_completed_
      -- 
    ra_1218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_615_inst_ack_0, ack => convTranspose_CP_34_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	475 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_update_completed_
      -- 
    ca_1223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_615_inst_ack_1, ack => convTranspose_CP_34_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	128 
    -- CP-element group 161: 	132 
    -- CP-element group 161: 	136 
    -- CP-element group 161: 	140 
    -- CP-element group 161: 	144 
    -- CP-element group 161: 	148 
    -- CP-element group 161: 	152 
    -- CP-element group 161: 	156 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/ptr_deref_623_Split/$exit
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/word_access_start/word_0/rr
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/word_access_start/word_0/$entry
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/word_access_start/$entry
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/ptr_deref_623_Split/split_ack
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/ptr_deref_623_Split/split_req
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/ptr_deref_623_Split/$entry
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_sample_start_
      -- 
    rr_1261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(161), ack => ptr_deref_623_store_0_req_0); -- 
    convTranspose_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(128) & convTranspose_CP_34_elements(132) & convTranspose_CP_34_elements(136) & convTranspose_CP_34_elements(140) & convTranspose_CP_34_elements(144) & convTranspose_CP_34_elements(148) & convTranspose_CP_34_elements(152) & convTranspose_CP_34_elements(156) & convTranspose_CP_34_elements(160);
      gj_convTranspose_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (5) 
      -- CP-element group 162: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/word_access_start/word_0/ra
      -- CP-element group 162: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/word_access_start/word_0/$exit
      -- CP-element group 162: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/word_access_start/$exit
      -- CP-element group 162: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_sample_completed_
      -- 
    ra_1262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_623_store_0_ack_0, ack => convTranspose_CP_34_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	475 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/word_access_complete/word_0/ca
      -- CP-element group 163: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/word_access_complete/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/word_access_complete/$exit
      -- CP-element group 163: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_update_completed_
      -- 
    ca_1273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_623_store_0_ack_1, ack => convTranspose_CP_34_elements(163)); -- 
    -- CP-element group 164:  branch  join  transition  place  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: 	125 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (10) 
      -- CP-element group 164: 	 branch_block_stmt_38/R_exitcond3_638_place
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637_if_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636__exit__
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637__entry__
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637_eval_test/branch_req
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637_eval_test/$exit
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637_eval_test/$entry
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637_dead_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_38/if_stmt_637_else_link/$entry
      -- CP-element group 164: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/$exit
      -- 
    branch_req_1281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(164), ack => if_stmt_637_branch_req_0); -- 
    convTranspose_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(163) & convTranspose_CP_34_elements(125);
      gj_convTranspose_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  merge  transition  place  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	469 
    -- CP-element group 165:  members (13) 
      -- CP-element group 165: 	 branch_block_stmt_38/merge_stmt_427__exit__
      -- CP-element group 165: 	 branch_block_stmt_38/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader
      -- CP-element group 165: 	 branch_block_stmt_38/if_stmt_637_if_link/if_choice_transition
      -- CP-element group 165: 	 branch_block_stmt_38/if_stmt_637_if_link/$exit
      -- CP-element group 165: 	 branch_block_stmt_38/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit
      -- CP-element group 165: 	 branch_block_stmt_38/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_38/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 165: 	 branch_block_stmt_38/merge_stmt_427_PhiReqMerge
      -- CP-element group 165: 	 branch_block_stmt_38/merge_stmt_427_PhiAck/$entry
      -- CP-element group 165: 	 branch_block_stmt_38/merge_stmt_427_PhiAck/$exit
      -- CP-element group 165: 	 branch_block_stmt_38/merge_stmt_427_PhiAck/dummy
      -- CP-element group 165: 	 branch_block_stmt_38/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 165: 	 branch_block_stmt_38/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_637_branch_ack_1, ack => convTranspose_CP_34_elements(165)); -- 
    -- CP-element group 166:  fork  transition  place  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	471 
    -- CP-element group 166: 	472 
    -- CP-element group 166:  members (12) 
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody
      -- CP-element group 166: 	 branch_block_stmt_38/if_stmt_637_else_link/else_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_38/if_stmt_637_else_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_637_branch_ack_0, ack => convTranspose_CP_34_elements(166)); -- 
    rr_3506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(166), ack => type_cast_480_inst_req_0); -- 
    cr_3511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(166), ack => type_cast_480_inst_req_1); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	121 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Sample/ra
      -- CP-element group 167: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_sample_completed_
      -- 
    ra_1304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_664_inst_ack_0, ack => convTranspose_CP_34_elements(167)); -- 
    -- CP-element group 168:  transition  place  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	121 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	476 
    -- CP-element group 168:  members (9) 
      -- CP-element group 168: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678__exit__
      -- CP-element group 168: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196
      -- CP-element group 168: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/type_cast_664_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_38/assign_stmt_649_to_assign_stmt_678/$exit
      -- CP-element group 168: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/$entry
      -- CP-element group 168: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_681/$entry
      -- CP-element group 168: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/$entry
      -- 
    ca_1309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_664_inst_ack_1, ack => convTranspose_CP_34_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	481 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	208 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Sample/ack
      -- CP-element group 169: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_sample_complete
      -- 
    ack_1338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_693_index_offset_ack_0, ack => convTranspose_CP_34_elements(169)); -- 
    -- CP-element group 170:  transition  input  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	481 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (11) 
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Update/ack
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_request/req
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_request/$entry
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_offset_calculated
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_base_plus_offset/sum_rename_ack
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_base_plus_offset/$entry
      -- 
    ack_1343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_693_index_offset_ack_1, ack => convTranspose_CP_34_elements(170)); -- 
    req_1352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(170), ack => addr_of_694_final_reg_req_0); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_request/$exit
      -- CP-element group 171: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_request/ack
      -- CP-element group 171: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_sample_completed_
      -- 
    ack_1353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_694_final_reg_ack_0, ack => convTranspose_CP_34_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	481 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	205 
    -- CP-element group 172:  members (19) 
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_complete/ack
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_complete/$exit
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_word_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_address_resized
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_addr_resize/$entry
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_addr_resize/$exit
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_addr_resize/base_resize_req
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_addr_resize/base_resize_ack
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_word_addrgen/$entry
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_word_addrgen/$exit
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_word_addrgen/root_register_req
      -- CP-element group 172: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_word_addrgen/root_register_ack
      -- 
    ack_1358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_694_final_reg_ack_1, ack => convTranspose_CP_34_elements(172)); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	481 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_update_start_
      -- CP-element group 173: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Update/cr
      -- CP-element group 173: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Sample/ra
      -- 
    ra_1367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_697_inst_ack_0, ack => convTranspose_CP_34_elements(173)); -- 
    cr_1371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(173), ack => RPIPE_ConvTranspose_input_pipe_697_inst_req_1); -- 
    -- CP-element group 174:  fork  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	177 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (9) 
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Update/ca
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Sample/$entry
      -- 
    ca_1372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_697_inst_ack_1, ack => convTranspose_CP_34_elements(174)); -- 
    rr_1394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(174), ack => RPIPE_ConvTranspose_input_pipe_710_inst_req_0); -- 
    rr_1380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(174), ack => type_cast_701_inst_req_0); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Sample/$exit
      -- 
    ra_1381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_701_inst_ack_0, ack => convTranspose_CP_34_elements(175)); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	481 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	205 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Update/$exit
      -- 
    ca_1386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_701_inst_ack_1, ack => convTranspose_CP_34_elements(176)); -- 
    -- CP-element group 177:  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	174 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_update_start_
      -- CP-element group 177: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_sample_completed_
      -- 
    ra_1395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_710_inst_ack_0, ack => convTranspose_CP_34_elements(177)); -- 
    cr_1399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(177), ack => RPIPE_ConvTranspose_input_pipe_710_inst_req_1); -- 
    -- CP-element group 178:  fork  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178: 	181 
    -- CP-element group 178:  members (9) 
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_710_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Sample/rr
      -- CP-element group 178: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Sample/$entry
      -- 
    ca_1400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_710_inst_ack_1, ack => convTranspose_CP_34_elements(178)); -- 
    rr_1408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(178), ack => type_cast_714_inst_req_0); -- 
    rr_1422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(178), ack => RPIPE_ConvTranspose_input_pipe_728_inst_req_0); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Sample/$exit
      -- 
    ra_1409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_714_inst_ack_0, ack => convTranspose_CP_34_elements(179)); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	481 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	205 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Update/$exit
      -- 
    ca_1414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_714_inst_ack_1, ack => convTranspose_CP_34_elements(180)); -- 
    -- CP-element group 181:  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	178 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (6) 
      -- CP-element group 181: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_update_start_
      -- CP-element group 181: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Update/cr
      -- CP-element group 181: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Sample/$exit
      -- 
    ra_1423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_728_inst_ack_0, ack => convTranspose_CP_34_elements(181)); -- 
    cr_1427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(181), ack => RPIPE_ConvTranspose_input_pipe_728_inst_req_1); -- 
    -- CP-element group 182:  fork  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182: 	185 
    -- CP-element group 182:  members (9) 
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Sample/rr
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_728_Update/$exit
      -- 
    ca_1428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_728_inst_ack_1, ack => convTranspose_CP_34_elements(182)); -- 
    rr_1436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(182), ack => type_cast_732_inst_req_0); -- 
    rr_1450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(182), ack => RPIPE_ConvTranspose_input_pipe_746_inst_req_0); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_sample_completed_
      -- 
    ra_1437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_732_inst_ack_0, ack => convTranspose_CP_34_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	481 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	205 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Update/$exit
      -- 
    ca_1442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_732_inst_ack_1, ack => convTranspose_CP_34_elements(184)); -- 
    -- CP-element group 185:  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	182 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Update/cr
      -- CP-element group 185: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_update_start_
      -- CP-element group 185: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_sample_completed_
      -- 
    ra_1451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_746_inst_ack_0, ack => convTranspose_CP_34_elements(185)); -- 
    cr_1455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(185), ack => RPIPE_ConvTranspose_input_pipe_746_inst_req_1); -- 
    -- CP-element group 186:  fork  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186: 	189 
    -- CP-element group 186:  members (9) 
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_746_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Sample/rr
      -- 
    ca_1456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_746_inst_ack_1, ack => convTranspose_CP_34_elements(186)); -- 
    rr_1464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(186), ack => type_cast_750_inst_req_0); -- 
    rr_1478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(186), ack => RPIPE_ConvTranspose_input_pipe_764_inst_req_0); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Sample/ra
      -- 
    ra_1465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_750_inst_ack_0, ack => convTranspose_CP_34_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	481 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	205 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Update/ca
      -- 
    ca_1470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_750_inst_ack_1, ack => convTranspose_CP_34_elements(188)); -- 
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	186 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_update_start_
      -- CP-element group 189: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Update/cr
      -- 
    ra_1479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_764_inst_ack_0, ack => convTranspose_CP_34_elements(189)); -- 
    cr_1483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(189), ack => RPIPE_ConvTranspose_input_pipe_764_inst_req_1); -- 
    -- CP-element group 190:  fork  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190: 	193 
    -- CP-element group 190:  members (9) 
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_764_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Sample/rr
      -- 
    ca_1484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_764_inst_ack_1, ack => convTranspose_CP_34_elements(190)); -- 
    rr_1492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(190), ack => type_cast_768_inst_req_0); -- 
    rr_1506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(190), ack => RPIPE_ConvTranspose_input_pipe_782_inst_req_0); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Sample/ra
      -- 
    ra_1493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_768_inst_ack_0, ack => convTranspose_CP_34_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	481 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	205 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Update/ca
      -- 
    ca_1498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_768_inst_ack_1, ack => convTranspose_CP_34_elements(192)); -- 
    -- CP-element group 193:  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	190 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (6) 
      -- CP-element group 193: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_update_start_
      -- CP-element group 193: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Update/$entry
      -- CP-element group 193: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Update/cr
      -- 
    ra_1507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_782_inst_ack_0, ack => convTranspose_CP_34_elements(193)); -- 
    cr_1511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(193), ack => RPIPE_ConvTranspose_input_pipe_782_inst_req_1); -- 
    -- CP-element group 194:  fork  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: 	197 
    -- CP-element group 194:  members (9) 
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_782_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Sample/rr
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Sample/rr
      -- 
    ca_1512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_782_inst_ack_1, ack => convTranspose_CP_34_elements(194)); -- 
    rr_1520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(194), ack => type_cast_786_inst_req_0); -- 
    rr_1534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(194), ack => RPIPE_ConvTranspose_input_pipe_800_inst_req_0); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Sample/ra
      -- 
    ra_1521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_786_inst_ack_0, ack => convTranspose_CP_34_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	481 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	205 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Update/ca
      -- 
    ca_1526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_786_inst_ack_1, ack => convTranspose_CP_34_elements(196)); -- 
    -- CP-element group 197:  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	194 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (6) 
      -- CP-element group 197: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_update_start_
      -- CP-element group 197: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Update/cr
      -- 
    ra_1535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_800_inst_ack_0, ack => convTranspose_CP_34_elements(197)); -- 
    cr_1539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(197), ack => RPIPE_ConvTranspose_input_pipe_800_inst_req_1); -- 
    -- CP-element group 198:  fork  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198: 	201 
    -- CP-element group 198:  members (9) 
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_800_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Sample/rr
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Sample/rr
      -- 
    ca_1540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_800_inst_ack_1, ack => convTranspose_CP_34_elements(198)); -- 
    rr_1548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(198), ack => type_cast_804_inst_req_0); -- 
    rr_1562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(198), ack => RPIPE_ConvTranspose_input_pipe_818_inst_req_0); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Sample/ra
      -- 
    ra_1549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_804_inst_ack_0, ack => convTranspose_CP_34_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	481 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	205 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Update/ca
      -- 
    ca_1554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_804_inst_ack_1, ack => convTranspose_CP_34_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	198 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_update_start_
      -- CP-element group 201: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Sample/ra
      -- CP-element group 201: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Update/cr
      -- 
    ra_1563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_818_inst_ack_0, ack => convTranspose_CP_34_elements(201)); -- 
    cr_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(201), ack => RPIPE_ConvTranspose_input_pipe_818_inst_req_1); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_818_Update/ca
      -- CP-element group 202: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Sample/rr
      -- 
    ca_1568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_818_inst_ack_1, ack => convTranspose_CP_34_elements(202)); -- 
    rr_1576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(202), ack => type_cast_822_inst_req_0); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Sample/ra
      -- 
    ra_1577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_822_inst_ack_0, ack => convTranspose_CP_34_elements(203)); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	481 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Update/ca
      -- 
    ca_1582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_822_inst_ack_1, ack => convTranspose_CP_34_elements(204)); -- 
    -- CP-element group 205:  join  transition  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	180 
    -- CP-element group 205: 	184 
    -- CP-element group 205: 	188 
    -- CP-element group 205: 	172 
    -- CP-element group 205: 	176 
    -- CP-element group 205: 	192 
    -- CP-element group 205: 	196 
    -- CP-element group 205: 	200 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (9) 
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/ptr_deref_830_Split/$entry
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/ptr_deref_830_Split/$exit
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/ptr_deref_830_Split/split_req
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/ptr_deref_830_Split/split_ack
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/word_access_start/$entry
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/word_access_start/word_0/$entry
      -- CP-element group 205: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/word_access_start/word_0/rr
      -- 
    rr_1620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(205), ack => ptr_deref_830_store_0_req_0); -- 
    convTranspose_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(180) & convTranspose_CP_34_elements(184) & convTranspose_CP_34_elements(188) & convTranspose_CP_34_elements(172) & convTranspose_CP_34_elements(176) & convTranspose_CP_34_elements(192) & convTranspose_CP_34_elements(196) & convTranspose_CP_34_elements(200) & convTranspose_CP_34_elements(204);
      gj_convTranspose_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (5) 
      -- CP-element group 206: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_sample_completed_
      -- CP-element group 206: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/word_access_start/$exit
      -- CP-element group 206: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/word_access_start/word_0/$exit
      -- CP-element group 206: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Sample/word_access_start/word_0/ra
      -- 
    ra_1621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_830_store_0_ack_0, ack => convTranspose_CP_34_elements(206)); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	481 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/word_access_complete/$exit
      -- CP-element group 207: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/word_access_complete/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/word_access_complete/word_0/ca
      -- 
    ca_1632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_830_store_0_ack_1, ack => convTranspose_CP_34_elements(207)); -- 
    -- CP-element group 208:  branch  join  transition  place  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: 	169 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (10) 
      -- CP-element group 208: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843__exit__
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844__entry__
      -- CP-element group 208: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/$exit
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844_dead_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844_eval_test/$entry
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844_eval_test/$exit
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844_eval_test/branch_req
      -- CP-element group 208: 	 branch_block_stmt_38/R_exitcond2_845_place
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844_if_link/$entry
      -- CP-element group 208: 	 branch_block_stmt_38/if_stmt_844_else_link/$entry
      -- 
    branch_req_1640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(208), ack => if_stmt_844_branch_req_0); -- 
    convTranspose_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(207) & convTranspose_CP_34_elements(169);
      gj_convTranspose_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  merge  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	482 
    -- CP-element group 209:  members (13) 
      -- CP-element group 209: 	 branch_block_stmt_38/merge_stmt_850__exit__
      -- CP-element group 209: 	 branch_block_stmt_38/forx_xend250x_xloopexit_forx_xend250
      -- CP-element group 209: 	 branch_block_stmt_38/if_stmt_844_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_38/if_stmt_844_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_38/forx_xbody196_forx_xend250x_xloopexit
      -- CP-element group 209: 	 branch_block_stmt_38/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_38/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_38/merge_stmt_850_PhiReqMerge
      -- CP-element group 209: 	 branch_block_stmt_38/merge_stmt_850_PhiAck/$entry
      -- CP-element group 209: 	 branch_block_stmt_38/merge_stmt_850_PhiAck/$exit
      -- CP-element group 209: 	 branch_block_stmt_38/merge_stmt_850_PhiAck/dummy
      -- CP-element group 209: 	 branch_block_stmt_38/forx_xend250x_xloopexit_forx_xend250_PhiReq/$entry
      -- CP-element group 209: 	 branch_block_stmt_38/forx_xend250x_xloopexit_forx_xend250_PhiReq/$exit
      -- 
    if_choice_transition_1645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_844_branch_ack_1, ack => convTranspose_CP_34_elements(209)); -- 
    -- CP-element group 210:  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	477 
    -- CP-element group 210: 	478 
    -- CP-element group 210:  members (12) 
      -- CP-element group 210: 	 branch_block_stmt_38/if_stmt_844_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_38/if_stmt_844_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_844_branch_ack_0, ack => convTranspose_CP_34_elements(210)); -- 
    rr_3560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(210), ack => type_cast_687_inst_req_0); -- 
    cr_3565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(210), ack => type_cast_687_inst_req_1); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	482 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Sample/ra
      -- 
    ra_1663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_855_inst_ack_0, ack => convTranspose_CP_34_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	482 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	217 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Update/ca
      -- 
    ca_1668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_855_inst_ack_1, ack => convTranspose_CP_34_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	482 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Sample/ra
      -- 
    ra_1677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_859_inst_ack_0, ack => convTranspose_CP_34_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	482 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	217 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Update/ca
      -- 
    ca_1682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_859_inst_ack_1, ack => convTranspose_CP_34_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	482 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Sample/ra
      -- 
    ra_1691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_863_inst_ack_0, ack => convTranspose_CP_34_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	482 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Update/ca
      -- 
    ca_1696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_863_inst_ack_1, ack => convTranspose_CP_34_elements(216)); -- 
    -- CP-element group 217:  branch  join  transition  place  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	212 
    -- CP-element group 217: 	214 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (10) 
      -- CP-element group 217: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880__exit__
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881__entry__
      -- CP-element group 217: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/$exit
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881_dead_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881_eval_test/$entry
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881_eval_test/$exit
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881_eval_test/branch_req
      -- CP-element group 217: 	 branch_block_stmt_38/R_cmp264505_882_place
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881_if_link/$entry
      -- CP-element group 217: 	 branch_block_stmt_38/if_stmt_881_else_link/$entry
      -- 
    branch_req_1704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(217), ack => if_stmt_881_branch_req_0); -- 
    convTranspose_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(212) & convTranspose_CP_34_elements(214) & convTranspose_CP_34_elements(216);
      gj_convTranspose_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: 	221 
    -- CP-element group 218:  members (18) 
      -- CP-element group 218: 	 branch_block_stmt_38/merge_stmt_887__exit__
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922__entry__
      -- CP-element group 218: 	 branch_block_stmt_38/if_stmt_881_if_link/$exit
      -- CP-element group 218: 	 branch_block_stmt_38/if_stmt_881_if_link/if_choice_transition
      -- CP-element group 218: 	 branch_block_stmt_38/forx_xend250_bbx_xnph507
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/$entry
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_update_start_
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Sample/rr
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Update/cr
      -- CP-element group 218: 	 branch_block_stmt_38/forx_xend250_bbx_xnph507_PhiReq/$entry
      -- CP-element group 218: 	 branch_block_stmt_38/forx_xend250_bbx_xnph507_PhiReq/$exit
      -- CP-element group 218: 	 branch_block_stmt_38/merge_stmt_887_PhiReqMerge
      -- CP-element group 218: 	 branch_block_stmt_38/merge_stmt_887_PhiAck/$entry
      -- CP-element group 218: 	 branch_block_stmt_38/merge_stmt_887_PhiAck/$exit
      -- CP-element group 218: 	 branch_block_stmt_38/merge_stmt_887_PhiAck/dummy
      -- 
    if_choice_transition_1709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_881_branch_ack_1, ack => convTranspose_CP_34_elements(218)); -- 
    rr_1726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(218), ack => type_cast_908_inst_req_0); -- 
    cr_1731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(218), ack => type_cast_908_inst_req_1); -- 
    -- CP-element group 219:  transition  place  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	489 
    -- CP-element group 219:  members (5) 
      -- CP-element group 219: 	 branch_block_stmt_38/if_stmt_881_else_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_38/if_stmt_881_else_link/else_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_38/forx_xend250_forx_xend273
      -- CP-element group 219: 	 branch_block_stmt_38/forx_xend250_forx_xend273_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_38/forx_xend250_forx_xend273_PhiReq/$exit
      -- 
    else_choice_transition_1713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_881_branch_ack_0, ack => convTranspose_CP_34_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Sample/ra
      -- 
    ra_1727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_908_inst_ack_0, ack => convTranspose_CP_34_elements(220)); -- 
    -- CP-element group 221:  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	218 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	483 
    -- CP-element group 221:  members (9) 
      -- CP-element group 221: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922__exit__
      -- CP-element group 221: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266
      -- CP-element group 221: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/$exit
      -- CP-element group 221: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_38/assign_stmt_893_to_assign_stmt_922/type_cast_908_Update/ca
      -- CP-element group 221: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_925/$entry
      -- CP-element group 221: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/$entry
      -- 
    ca_1732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_908_inst_ack_1, ack => convTranspose_CP_34_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	488 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	228 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_sample_complete
      -- CP-element group 222: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Sample/ack
      -- 
    ack_1761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_937_index_offset_ack_0, ack => convTranspose_CP_34_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	488 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (11) 
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_root_address_calculated
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_offset_calculated
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Update/ack
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_base_plus_offset/$entry
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_base_plus_offset/$exit
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_base_plus_offset/sum_rename_req
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_base_plus_offset/sum_rename_ack
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_request/$entry
      -- CP-element group 223: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_request/req
      -- 
    ack_1766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_937_index_offset_ack_1, ack => convTranspose_CP_34_elements(223)); -- 
    req_1775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(223), ack => addr_of_938_final_reg_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_request/$exit
      -- CP-element group 224: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_request/ack
      -- 
    ack_1776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_938_final_reg_ack_0, ack => convTranspose_CP_34_elements(224)); -- 
    -- CP-element group 225:  join  fork  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	488 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (28) 
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_complete/$exit
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_complete/ack
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_word_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_address_resized
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_addr_resize/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_addr_resize/$exit
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_addr_resize/base_resize_req
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_addr_resize/base_resize_ack
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_plus_offset/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_word_addrgen/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_word_addrgen/$exit
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_word_addrgen/root_register_req
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_word_addrgen/root_register_ack
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/ptr_deref_941_Split/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/ptr_deref_941_Split/$exit
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/ptr_deref_941_Split/split_req
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/ptr_deref_941_Split/split_ack
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/word_access_start/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/word_access_start/word_0/$entry
      -- CP-element group 225: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/word_access_start/word_0/rr
      -- 
    ack_1781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_938_final_reg_ack_1, ack => convTranspose_CP_34_elements(225)); -- 
    rr_1819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(225), ack => ptr_deref_941_store_0_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/word_access_start/$exit
      -- CP-element group 226: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/word_access_start/word_0/$exit
      -- CP-element group 226: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Sample/word_access_start/word_0/ra
      -- 
    ra_1820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_941_store_0_ack_0, ack => convTranspose_CP_34_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	488 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/word_access_complete/$exit
      -- CP-element group 227: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/word_access_complete/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/word_access_complete/word_0/ca
      -- 
    ca_1831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_941_store_0_ack_1, ack => convTranspose_CP_34_elements(227)); -- 
    -- CP-element group 228:  branch  join  transition  place  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	222 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (10) 
      -- CP-element group 228: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955__exit__
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956__entry__
      -- CP-element group 228: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/$exit
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956_dead_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956_eval_test/$entry
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956_eval_test/$exit
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956_eval_test/branch_req
      -- CP-element group 228: 	 branch_block_stmt_38/R_exitcond_957_place
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956_if_link/$entry
      -- CP-element group 228: 	 branch_block_stmt_38/if_stmt_956_else_link/$entry
      -- 
    branch_req_1839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(228), ack => if_stmt_956_branch_req_0); -- 
    convTranspose_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(222) & convTranspose_CP_34_elements(227);
      gj_convTranspose_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  merge  transition  place  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	489 
    -- CP-element group 229:  members (13) 
      -- CP-element group 229: 	 branch_block_stmt_38/merge_stmt_962__exit__
      -- CP-element group 229: 	 branch_block_stmt_38/forx_xend273x_xloopexit_forx_xend273
      -- CP-element group 229: 	 branch_block_stmt_38/if_stmt_956_if_link/$exit
      -- CP-element group 229: 	 branch_block_stmt_38/if_stmt_956_if_link/if_choice_transition
      -- CP-element group 229: 	 branch_block_stmt_38/forx_xbody266_forx_xend273x_xloopexit
      -- CP-element group 229: 	 branch_block_stmt_38/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_38/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$exit
      -- CP-element group 229: 	 branch_block_stmt_38/merge_stmt_962_PhiReqMerge
      -- CP-element group 229: 	 branch_block_stmt_38/merge_stmt_962_PhiAck/$entry
      -- CP-element group 229: 	 branch_block_stmt_38/merge_stmt_962_PhiAck/$exit
      -- CP-element group 229: 	 branch_block_stmt_38/merge_stmt_962_PhiAck/dummy
      -- CP-element group 229: 	 branch_block_stmt_38/forx_xend273x_xloopexit_forx_xend273_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_38/forx_xend273x_xloopexit_forx_xend273_PhiReq/$exit
      -- 
    if_choice_transition_1844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_956_branch_ack_1, ack => convTranspose_CP_34_elements(229)); -- 
    -- CP-element group 230:  fork  transition  place  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	484 
    -- CP-element group 230: 	485 
    -- CP-element group 230:  members (12) 
      -- CP-element group 230: 	 branch_block_stmt_38/if_stmt_956_else_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_38/if_stmt_956_else_link/else_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_956_branch_ack_0, ack => convTranspose_CP_34_elements(230)); -- 
    rr_3637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(230), ack => type_cast_928_inst_req_0); -- 
    cr_3642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(230), ack => type_cast_928_inst_req_1); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	489 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Sample/cra
      -- 
    cra_1862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_967_call_ack_0, ack => convTranspose_CP_34_elements(231)); -- 
    -- CP-element group 232:  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	489 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Update/cca
      -- CP-element group 232: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Sample/rr
      -- 
    cca_1867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_967_call_ack_1, ack => convTranspose_CP_34_elements(232)); -- 
    rr_1875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(232), ack => type_cast_972_inst_req_0); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Sample/ra
      -- 
    ra_1876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_972_inst_ack_0, ack => convTranspose_CP_34_elements(233)); -- 
    -- CP-element group 234:  fork  transition  place  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	489 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	263 
    -- CP-element group 234: 	281 
    -- CP-element group 234: 	282 
    -- CP-element group 234: 	286 
    -- CP-element group 234: 	287 
    -- CP-element group 234: 	297 
    -- CP-element group 234: 	315 
    -- CP-element group 234: 	316 
    -- CP-element group 234: 	320 
    -- CP-element group 234: 	321 
    -- CP-element group 234: 	331 
    -- CP-element group 234: 	349 
    -- CP-element group 234: 	350 
    -- CP-element group 234: 	354 
    -- CP-element group 234: 	355 
    -- CP-element group 234: 	365 
    -- CP-element group 234: 	367 
    -- CP-element group 234: 	369 
    -- CP-element group 234: 	371 
    -- CP-element group 234: 	235 
    -- CP-element group 234:  members (67) 
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1019_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973__exit__
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198__entry__
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1061_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1075_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1019_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1075_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1019_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1075_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1054_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1054_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1054_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1054_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1054_update_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1054_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1061_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1061_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1061_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1061_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1061_update_start_
      -- CP-element group 234: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/$exit
      -- CP-element group 234: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Update/ca
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_975_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_975_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_975_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1110_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1110_update_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1110_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1110_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1110_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1110_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1117_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1117_update_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1117_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1117_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1117_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1117_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1131_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1131_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1131_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1166_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1166_update_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1166_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1166_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1166_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1166_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1173_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1173_update_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1173_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1173_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1173_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1173_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block0_done_1188_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block0_done_1188_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block0_done_1188_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block1_done_1191_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block1_done_1191_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block1_done_1191_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block2_done_1194_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block2_done_1194_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block2_done_1194_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block3_done_1197_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block3_done_1197_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block3_done_1197_Sample/rr
      -- 
    ca_1881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_972_inst_ack_1, ack => convTranspose_CP_34_elements(234)); -- 
    req_2312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => WPIPE_Block2_start_1075_inst_req_0); -- 
    req_2088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => WPIPE_Block1_start_1019_inst_req_0); -- 
    cr_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1054_inst_req_1); -- 
    rr_2214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1054_inst_req_0); -- 
    cr_2247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1061_inst_req_1); -- 
    rr_2242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1061_inst_req_0); -- 
    req_1892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => WPIPE_Block0_start_975_inst_req_0); -- 
    rr_2438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1110_inst_req_0); -- 
    cr_2443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1110_inst_req_1); -- 
    rr_2466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1117_inst_req_0); -- 
    cr_2471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1117_inst_req_1); -- 
    req_2536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => WPIPE_Block3_start_1131_inst_req_0); -- 
    rr_2662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1166_inst_req_0); -- 
    cr_2667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1166_inst_req_1); -- 
    rr_2690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1173_inst_req_0); -- 
    cr_2695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => type_cast_1173_inst_req_1); -- 
    rr_2760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => RPIPE_Block0_done_1188_inst_req_0); -- 
    rr_2774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => RPIPE_Block1_done_1191_inst_req_0); -- 
    rr_2788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => RPIPE_Block2_done_1194_inst_req_0); -- 
    rr_2802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(234), ack => RPIPE_Block3_done_1197_inst_req_0); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_975_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_975_update_start_
      -- CP-element group 235: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_975_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_975_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_975_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_975_Update/req
      -- 
    ack_1893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_975_inst_ack_0, ack => convTranspose_CP_34_elements(235)); -- 
    req_1897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(235), ack => WPIPE_Block0_start_975_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_978_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_978_Sample/req
      -- CP-element group 236: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_975_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_975_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_975_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_978_sample_start_
      -- 
    ack_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_975_inst_ack_1, ack => convTranspose_CP_34_elements(236)); -- 
    req_1906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(236), ack => WPIPE_Block0_start_978_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_978_Update/req
      -- CP-element group 237: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_978_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_978_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_978_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_978_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_978_update_start_
      -- 
    ack_1907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_978_inst_ack_0, ack => convTranspose_CP_34_elements(237)); -- 
    req_1911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(237), ack => WPIPE_Block0_start_978_inst_req_1); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_978_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_978_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_981_Sample/req
      -- CP-element group 238: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_981_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_981_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_978_update_completed_
      -- 
    ack_1912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_978_inst_ack_1, ack => convTranspose_CP_34_elements(238)); -- 
    req_1920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(238), ack => WPIPE_Block0_start_981_inst_req_0); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_981_update_start_
      -- CP-element group 239: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_981_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_981_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_981_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_981_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_981_Update/req
      -- 
    ack_1921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_981_inst_ack_0, ack => convTranspose_CP_34_elements(239)); -- 
    req_1925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(239), ack => WPIPE_Block0_start_981_inst_req_1); -- 
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_981_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_981_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_981_Update/ack
      -- CP-element group 240: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_984_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_984_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_984_Sample/req
      -- 
    ack_1926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_981_inst_ack_1, ack => convTranspose_CP_34_elements(240)); -- 
    req_1934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(240), ack => WPIPE_Block0_start_984_inst_req_0); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_984_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_984_update_start_
      -- CP-element group 241: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_984_Update/req
      -- CP-element group 241: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_984_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_984_Sample/ack
      -- CP-element group 241: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_984_Sample/$exit
      -- 
    ack_1935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_984_inst_ack_0, ack => convTranspose_CP_34_elements(241)); -- 
    req_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(241), ack => WPIPE_Block0_start_984_inst_req_1); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_984_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_987_Sample/req
      -- CP-element group 242: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_987_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_987_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_984_Update/ack
      -- CP-element group 242: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_984_Update/$exit
      -- 
    ack_1940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_984_inst_ack_1, ack => convTranspose_CP_34_elements(242)); -- 
    req_1948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(242), ack => WPIPE_Block0_start_987_inst_req_0); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_987_Update/req
      -- CP-element group 243: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_987_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_987_Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_987_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_987_update_start_
      -- CP-element group 243: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_987_sample_completed_
      -- 
    ack_1949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_987_inst_ack_0, ack => convTranspose_CP_34_elements(243)); -- 
    req_1953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(243), ack => WPIPE_Block0_start_987_inst_req_1); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_987_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_990_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_987_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_990_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_990_Sample/req
      -- CP-element group 244: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_987_update_completed_
      -- 
    ack_1954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_987_inst_ack_1, ack => convTranspose_CP_34_elements(244)); -- 
    req_1962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(244), ack => WPIPE_Block0_start_990_inst_req_0); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_990_update_start_
      -- CP-element group 245: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_990_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_990_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_990_Sample/ack
      -- CP-element group 245: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_990_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_990_Update/req
      -- 
    ack_1963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_990_inst_ack_0, ack => convTranspose_CP_34_elements(245)); -- 
    req_1967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(245), ack => WPIPE_Block0_start_990_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_990_update_completed_
      -- CP-element group 246: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_990_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_993_Sample/req
      -- CP-element group 246: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_993_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_993_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_990_Update/ack
      -- 
    ack_1968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_990_inst_ack_1, ack => convTranspose_CP_34_elements(246)); -- 
    req_1976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(246), ack => WPIPE_Block0_start_993_inst_req_0); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_993_Update/req
      -- CP-element group 247: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_993_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_993_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_993_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_993_update_start_
      -- CP-element group 247: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_993_sample_completed_
      -- 
    ack_1977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_993_inst_ack_0, ack => convTranspose_CP_34_elements(247)); -- 
    req_1981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(247), ack => WPIPE_Block0_start_993_inst_req_1); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_993_Update/ack
      -- CP-element group 248: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_996_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_996_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_996_Sample/req
      -- CP-element group 248: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_993_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_993_update_completed_
      -- 
    ack_1982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_993_inst_ack_1, ack => convTranspose_CP_34_elements(248)); -- 
    req_1990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(248), ack => WPIPE_Block0_start_996_inst_req_0); -- 
    -- CP-element group 249:  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (6) 
      -- CP-element group 249: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_996_sample_completed_
      -- CP-element group 249: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_996_Sample/ack
      -- CP-element group 249: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_996_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_996_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_996_update_start_
      -- CP-element group 249: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_996_Update/req
      -- 
    ack_1991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_996_inst_ack_0, ack => convTranspose_CP_34_elements(249)); -- 
    req_1995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(249), ack => WPIPE_Block0_start_996_inst_req_1); -- 
    -- CP-element group 250:  transition  input  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (6) 
      -- CP-element group 250: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_996_update_completed_
      -- CP-element group 250: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_996_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_999_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_996_Update/ack
      -- CP-element group 250: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_999_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_999_Sample/req
      -- 
    ack_1996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_996_inst_ack_1, ack => convTranspose_CP_34_elements(250)); -- 
    req_2004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(250), ack => WPIPE_Block0_start_999_inst_req_0); -- 
    -- CP-element group 251:  transition  input  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_999_update_start_
      -- CP-element group 251: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_999_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_999_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_999_Sample/ack
      -- CP-element group 251: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_999_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_999_Update/req
      -- 
    ack_2005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_999_inst_ack_0, ack => convTranspose_CP_34_elements(251)); -- 
    req_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(251), ack => WPIPE_Block0_start_999_inst_req_1); -- 
    -- CP-element group 252:  transition  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (6) 
      -- CP-element group 252: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_999_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_999_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_999_Update/ack
      -- CP-element group 252: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1002_Sample/req
      -- CP-element group 252: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1002_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1002_sample_start_
      -- 
    ack_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_999_inst_ack_1, ack => convTranspose_CP_34_elements(252)); -- 
    req_2018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(252), ack => WPIPE_Block0_start_1002_inst_req_0); -- 
    -- CP-element group 253:  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1002_Update/req
      -- CP-element group 253: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1002_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1002_Sample/ack
      -- CP-element group 253: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1002_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1002_update_start_
      -- CP-element group 253: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1002_sample_completed_
      -- 
    ack_2019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1002_inst_ack_0, ack => convTranspose_CP_34_elements(253)); -- 
    req_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(253), ack => WPIPE_Block0_start_1002_inst_req_1); -- 
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (6) 
      -- CP-element group 254: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1006_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1002_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1002_Update/ack
      -- CP-element group 254: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1006_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1006_Sample/req
      -- CP-element group 254: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1002_update_completed_
      -- 
    ack_2024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1002_inst_ack_1, ack => convTranspose_CP_34_elements(254)); -- 
    req_2032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(254), ack => WPIPE_Block0_start_1006_inst_req_0); -- 
    -- CP-element group 255:  transition  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (6) 
      -- CP-element group 255: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1006_update_start_
      -- CP-element group 255: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1006_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1006_Update/req
      -- CP-element group 255: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1006_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1006_Sample/ack
      -- CP-element group 255: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1006_Update/$entry
      -- 
    ack_2033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1006_inst_ack_0, ack => convTranspose_CP_34_elements(255)); -- 
    req_2037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(255), ack => WPIPE_Block0_start_1006_inst_req_1); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1006_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1006_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1010_Sample/req
      -- CP-element group 256: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1010_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1010_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1006_Update/ack
      -- 
    ack_2038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1006_inst_ack_1, ack => convTranspose_CP_34_elements(256)); -- 
    req_2046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(256), ack => WPIPE_Block0_start_1010_inst_req_0); -- 
    -- CP-element group 257:  transition  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (6) 
      -- CP-element group 257: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1010_Update/req
      -- CP-element group 257: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1010_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1010_Sample/ack
      -- CP-element group 257: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1010_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1010_update_start_
      -- CP-element group 257: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1010_sample_completed_
      -- 
    ack_2047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1010_inst_ack_0, ack => convTranspose_CP_34_elements(257)); -- 
    req_2051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(257), ack => WPIPE_Block0_start_1010_inst_req_1); -- 
    -- CP-element group 258:  transition  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (6) 
      -- CP-element group 258: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1013_Sample/req
      -- CP-element group 258: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1013_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1013_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1010_Update/ack
      -- CP-element group 258: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1010_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1010_update_completed_
      -- 
    ack_2052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1010_inst_ack_1, ack => convTranspose_CP_34_elements(258)); -- 
    req_2060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(258), ack => WPIPE_Block0_start_1013_inst_req_0); -- 
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1013_Update/req
      -- CP-element group 259: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1013_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1013_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1013_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1013_update_start_
      -- CP-element group 259: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1013_sample_completed_
      -- 
    ack_2061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1013_inst_ack_0, ack => convTranspose_CP_34_elements(259)); -- 
    req_2065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(259), ack => WPIPE_Block0_start_1013_inst_req_1); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1016_Sample/req
      -- CP-element group 260: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1016_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1016_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1013_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1013_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1013_update_completed_
      -- 
    ack_2066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1013_inst_ack_1, ack => convTranspose_CP_34_elements(260)); -- 
    req_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(260), ack => WPIPE_Block0_start_1016_inst_req_0); -- 
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1016_Update/req
      -- CP-element group 261: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1016_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1016_Sample/ack
      -- CP-element group 261: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1016_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1016_update_start_
      -- CP-element group 261: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1016_sample_completed_
      -- 
    ack_2075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1016_inst_ack_0, ack => convTranspose_CP_34_elements(261)); -- 
    req_2079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(261), ack => WPIPE_Block0_start_1016_inst_req_1); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	373 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1016_Update/ack
      -- CP-element group 262: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1016_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block0_start_1016_update_completed_
      -- 
    ack_2080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1016_inst_ack_1, ack => convTranspose_CP_34_elements(262)); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	234 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1019_Update/req
      -- CP-element group 263: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1019_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1019_update_start_
      -- CP-element group 263: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1019_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1019_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1019_Sample/ack
      -- 
    ack_2089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1019_inst_ack_0, ack => convTranspose_CP_34_elements(263)); -- 
    req_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(263), ack => WPIPE_Block1_start_1019_inst_req_1); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1019_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1019_Update/ack
      -- CP-element group 264: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1022_Sample/req
      -- CP-element group 264: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1022_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1019_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1022_Sample/$entry
      -- 
    ack_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1019_inst_ack_1, ack => convTranspose_CP_34_elements(264)); -- 
    req_2102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(264), ack => WPIPE_Block1_start_1022_inst_req_0); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (6) 
      -- CP-element group 265: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1022_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1022_Update/$entry
      -- CP-element group 265: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1022_Sample/ack
      -- CP-element group 265: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1022_sample_completed_
      -- CP-element group 265: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1022_Update/req
      -- CP-element group 265: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1022_update_start_
      -- 
    ack_2103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1022_inst_ack_0, ack => convTranspose_CP_34_elements(265)); -- 
    req_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(265), ack => WPIPE_Block1_start_1022_inst_req_1); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1022_update_completed_
      -- CP-element group 266: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1022_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1022_Update/ack
      -- CP-element group 266: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1025_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1025_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1025_Sample/req
      -- 
    ack_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1022_inst_ack_1, ack => convTranspose_CP_34_elements(266)); -- 
    req_2116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(266), ack => WPIPE_Block1_start_1025_inst_req_0); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1025_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1025_update_start_
      -- CP-element group 267: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1025_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1025_Sample/ack
      -- CP-element group 267: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1025_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1025_Update/req
      -- 
    ack_2117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1025_inst_ack_0, ack => convTranspose_CP_34_elements(267)); -- 
    req_2121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(267), ack => WPIPE_Block1_start_1025_inst_req_1); -- 
    -- CP-element group 268:  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (6) 
      -- CP-element group 268: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1025_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1028_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1025_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1025_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1028_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1028_Sample/req
      -- 
    ack_2122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1025_inst_ack_1, ack => convTranspose_CP_34_elements(268)); -- 
    req_2130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(268), ack => WPIPE_Block1_start_1028_inst_req_0); -- 
    -- CP-element group 269:  transition  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (6) 
      -- CP-element group 269: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1028_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1028_sample_completed_
      -- CP-element group 269: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1028_update_start_
      -- CP-element group 269: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1028_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1028_Sample/ack
      -- CP-element group 269: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1028_Update/req
      -- 
    ack_2131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1028_inst_ack_0, ack => convTranspose_CP_34_elements(269)); -- 
    req_2135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(269), ack => WPIPE_Block1_start_1028_inst_req_1); -- 
    -- CP-element group 270:  transition  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1028_update_completed_
      -- CP-element group 270: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1031_Sample/req
      -- CP-element group 270: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1031_Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1031_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1028_Update/ack
      -- CP-element group 270: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1028_Update/$exit
      -- 
    ack_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1028_inst_ack_1, ack => convTranspose_CP_34_elements(270)); -- 
    req_2144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(270), ack => WPIPE_Block1_start_1031_inst_req_0); -- 
    -- CP-element group 271:  transition  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (6) 
      -- CP-element group 271: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1031_Update/req
      -- CP-element group 271: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1031_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1031_Sample/ack
      -- CP-element group 271: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1031_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1031_update_start_
      -- CP-element group 271: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1031_sample_completed_
      -- 
    ack_2145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1031_inst_ack_0, ack => convTranspose_CP_34_elements(271)); -- 
    req_2149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(271), ack => WPIPE_Block1_start_1031_inst_req_1); -- 
    -- CP-element group 272:  transition  input  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (6) 
      -- CP-element group 272: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1034_Sample/req
      -- CP-element group 272: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1034_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1034_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1031_Update/ack
      -- CP-element group 272: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1031_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1031_update_completed_
      -- 
    ack_2150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1031_inst_ack_1, ack => convTranspose_CP_34_elements(272)); -- 
    req_2158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(272), ack => WPIPE_Block1_start_1034_inst_req_0); -- 
    -- CP-element group 273:  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1034_Update/req
      -- CP-element group 273: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1034_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1034_Sample/ack
      -- CP-element group 273: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1034_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1034_update_start_
      -- CP-element group 273: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1034_sample_completed_
      -- 
    ack_2159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1034_inst_ack_0, ack => convTranspose_CP_34_elements(273)); -- 
    req_2163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(273), ack => WPIPE_Block1_start_1034_inst_req_1); -- 
    -- CP-element group 274:  transition  input  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (6) 
      -- CP-element group 274: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1037_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1037_Sample/req
      -- CP-element group 274: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1034_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1034_Update/ack
      -- CP-element group 274: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1037_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1034_update_completed_
      -- 
    ack_2164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1034_inst_ack_1, ack => convTranspose_CP_34_elements(274)); -- 
    req_2172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(274), ack => WPIPE_Block1_start_1037_inst_req_0); -- 
    -- CP-element group 275:  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1037_update_start_
      -- CP-element group 275: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1037_sample_completed_
      -- CP-element group 275: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1037_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1037_Update/req
      -- CP-element group 275: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1037_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1037_Sample/ack
      -- 
    ack_2173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1037_inst_ack_0, ack => convTranspose_CP_34_elements(275)); -- 
    req_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(275), ack => WPIPE_Block1_start_1037_inst_req_1); -- 
    -- CP-element group 276:  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1037_update_completed_
      -- CP-element group 276: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1040_Sample/req
      -- CP-element group 276: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1040_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1040_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1037_Update/ack
      -- CP-element group 276: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1037_Update/$exit
      -- 
    ack_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1037_inst_ack_1, ack => convTranspose_CP_34_elements(276)); -- 
    req_2186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(276), ack => WPIPE_Block1_start_1040_inst_req_0); -- 
    -- CP-element group 277:  transition  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1040_Update/req
      -- CP-element group 277: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1040_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1040_Sample/ack
      -- CP-element group 277: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1040_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1040_update_start_
      -- CP-element group 277: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1040_sample_completed_
      -- 
    ack_2187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1040_inst_ack_0, ack => convTranspose_CP_34_elements(277)); -- 
    req_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(277), ack => WPIPE_Block1_start_1040_inst_req_1); -- 
    -- CP-element group 278:  transition  input  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (6) 
      -- CP-element group 278: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1043_Sample/req
      -- CP-element group 278: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1043_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1043_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1040_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1040_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1040_update_completed_
      -- 
    ack_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1040_inst_ack_1, ack => convTranspose_CP_34_elements(278)); -- 
    req_2200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(278), ack => WPIPE_Block1_start_1043_inst_req_0); -- 
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1043_Update/req
      -- CP-element group 279: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1043_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1043_Sample/ack
      -- CP-element group 279: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1043_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1043_update_start_
      -- CP-element group 279: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1043_sample_completed_
      -- 
    ack_2201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1043_inst_ack_0, ack => convTranspose_CP_34_elements(279)); -- 
    req_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(279), ack => WPIPE_Block1_start_1043_inst_req_1); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	283 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1043_Update/ack
      -- CP-element group 280: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1043_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1043_update_completed_
      -- 
    ack_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1043_inst_ack_1, ack => convTranspose_CP_34_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	234 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1054_Sample/ra
      -- CP-element group 281: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1054_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1054_sample_completed_
      -- 
    ra_2215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1054_inst_ack_0, ack => convTranspose_CP_34_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	234 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1054_Update/ca
      -- CP-element group 282: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1054_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1054_update_completed_
      -- 
    ca_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1054_inst_ack_1, ack => convTranspose_CP_34_elements(282)); -- 
    -- CP-element group 283:  join  transition  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	280 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1056_Sample/req
      -- CP-element group 283: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1056_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1056_sample_start_
      -- 
    req_2228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(283), ack => WPIPE_Block1_start_1056_inst_req_0); -- 
    convTranspose_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(280) & convTranspose_CP_34_elements(282);
      gj_convTranspose_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  transition  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1056_sample_completed_
      -- CP-element group 284: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1056_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1056_update_start_
      -- CP-element group 284: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1056_Sample/ack
      -- CP-element group 284: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1056_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1056_Update/req
      -- 
    ack_2229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1056_inst_ack_0, ack => convTranspose_CP_34_elements(284)); -- 
    req_2233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(284), ack => WPIPE_Block1_start_1056_inst_req_1); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	288 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1056_update_completed_
      -- CP-element group 285: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1056_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1056_Update/ack
      -- 
    ack_2234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1056_inst_ack_1, ack => convTranspose_CP_34_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	234 
    -- CP-element group 286: successors 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1061_Sample/ra
      -- CP-element group 286: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1061_Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1061_sample_completed_
      -- 
    ra_2243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1061_inst_ack_0, ack => convTranspose_CP_34_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	234 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1061_Update/ca
      -- CP-element group 287: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1061_Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1061_update_completed_
      -- 
    ca_2248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1061_inst_ack_1, ack => convTranspose_CP_34_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	285 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1063_Sample/req
      -- CP-element group 288: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1063_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1063_sample_start_
      -- 
    req_2256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(288), ack => WPIPE_Block1_start_1063_inst_req_0); -- 
    convTranspose_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(285) & convTranspose_CP_34_elements(287);
      gj_convTranspose_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  transition  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (6) 
      -- CP-element group 289: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1063_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1063_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1063_Update/req
      -- CP-element group 289: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1063_Sample/ack
      -- CP-element group 289: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1063_update_start_
      -- CP-element group 289: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1063_sample_completed_
      -- 
    ack_2257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1063_inst_ack_0, ack => convTranspose_CP_34_elements(289)); -- 
    req_2261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(289), ack => WPIPE_Block1_start_1063_inst_req_1); -- 
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1063_Update/ack
      -- CP-element group 290: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1063_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1066_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1063_update_completed_
      -- CP-element group 290: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1066_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1066_Sample/$entry
      -- 
    ack_2262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1063_inst_ack_1, ack => convTranspose_CP_34_elements(290)); -- 
    req_2270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(290), ack => WPIPE_Block1_start_1066_inst_req_0); -- 
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1066_sample_completed_
      -- CP-element group 291: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1066_update_start_
      -- CP-element group 291: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1066_Update/req
      -- CP-element group 291: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1066_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1066_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1066_Sample/$exit
      -- 
    ack_2271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1066_inst_ack_0, ack => convTranspose_CP_34_elements(291)); -- 
    req_2275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(291), ack => WPIPE_Block1_start_1066_inst_req_1); -- 
    -- CP-element group 292:  transition  input  output  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (6) 
      -- CP-element group 292: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1069_sample_start_
      -- CP-element group 292: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1069_Sample/$entry
      -- CP-element group 292: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1066_Update/ack
      -- CP-element group 292: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1066_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1069_Sample/req
      -- CP-element group 292: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1066_update_completed_
      -- 
    ack_2276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1066_inst_ack_1, ack => convTranspose_CP_34_elements(292)); -- 
    req_2284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(292), ack => WPIPE_Block1_start_1069_inst_req_0); -- 
    -- CP-element group 293:  transition  input  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1069_Update/req
      -- CP-element group 293: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1069_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1069_sample_completed_
      -- CP-element group 293: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1069_update_start_
      -- CP-element group 293: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1069_Update/$entry
      -- CP-element group 293: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1069_Sample/ack
      -- 
    ack_2285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1069_inst_ack_0, ack => convTranspose_CP_34_elements(293)); -- 
    req_2289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(293), ack => WPIPE_Block1_start_1069_inst_req_1); -- 
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1069_Update/ack
      -- CP-element group 294: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1069_update_completed_
      -- CP-element group 294: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1069_Update/$exit
      -- CP-element group 294: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1072_Sample/req
      -- CP-element group 294: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1072_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1072_sample_start_
      -- 
    ack_2290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1069_inst_ack_1, ack => convTranspose_CP_34_elements(294)); -- 
    req_2298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(294), ack => WPIPE_Block1_start_1072_inst_req_0); -- 
    -- CP-element group 295:  transition  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (6) 
      -- CP-element group 295: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1072_Update/req
      -- CP-element group 295: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1072_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1072_Sample/ack
      -- CP-element group 295: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1072_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1072_update_start_
      -- CP-element group 295: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1072_sample_completed_
      -- 
    ack_2299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1072_inst_ack_0, ack => convTranspose_CP_34_elements(295)); -- 
    req_2303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(295), ack => WPIPE_Block1_start_1072_inst_req_1); -- 
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	373 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1072_Update/ack
      -- CP-element group 296: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1072_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block1_start_1072_update_completed_
      -- 
    ack_2304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1072_inst_ack_1, ack => convTranspose_CP_34_elements(296)); -- 
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	234 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1075_update_start_
      -- CP-element group 297: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1075_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1075_sample_completed_
      -- CP-element group 297: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1075_Update/req
      -- CP-element group 297: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1075_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1075_Sample/ack
      -- 
    ack_2313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1075_inst_ack_0, ack => convTranspose_CP_34_elements(297)); -- 
    req_2317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(297), ack => WPIPE_Block2_start_1075_inst_req_1); -- 
    -- CP-element group 298:  transition  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (6) 
      -- CP-element group 298: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1075_update_completed_
      -- CP-element group 298: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1078_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1075_Update/ack
      -- CP-element group 298: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1075_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1078_Sample/req
      -- CP-element group 298: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1078_Sample/$entry
      -- 
    ack_2318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1075_inst_ack_1, ack => convTranspose_CP_34_elements(298)); -- 
    req_2326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(298), ack => WPIPE_Block2_start_1078_inst_req_0); -- 
    -- CP-element group 299:  transition  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1078_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1078_Update/req
      -- CP-element group 299: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1078_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1078_Sample/ack
      -- CP-element group 299: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1078_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1078_update_start_
      -- 
    ack_2327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1078_inst_ack_0, ack => convTranspose_CP_34_elements(299)); -- 
    req_2331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(299), ack => WPIPE_Block2_start_1078_inst_req_1); -- 
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1081_sample_start_
      -- CP-element group 300: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1078_Update/ack
      -- CP-element group 300: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1078_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1081_Sample/req
      -- CP-element group 300: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1081_Sample/$entry
      -- CP-element group 300: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1078_update_completed_
      -- 
    ack_2332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1078_inst_ack_1, ack => convTranspose_CP_34_elements(300)); -- 
    req_2340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(300), ack => WPIPE_Block2_start_1081_inst_req_0); -- 
    -- CP-element group 301:  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (6) 
      -- CP-element group 301: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1081_sample_completed_
      -- CP-element group 301: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1081_Update/req
      -- CP-element group 301: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1081_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1081_Sample/ack
      -- CP-element group 301: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1081_Sample/$exit
      -- CP-element group 301: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1081_update_start_
      -- 
    ack_2341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1081_inst_ack_0, ack => convTranspose_CP_34_elements(301)); -- 
    req_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(301), ack => WPIPE_Block2_start_1081_inst_req_1); -- 
    -- CP-element group 302:  transition  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (6) 
      -- CP-element group 302: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1084_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1084_Sample/req
      -- CP-element group 302: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1081_Update/ack
      -- CP-element group 302: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1084_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1081_Update/$exit
      -- CP-element group 302: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1081_update_completed_
      -- 
    ack_2346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1081_inst_ack_1, ack => convTranspose_CP_34_elements(302)); -- 
    req_2354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(302), ack => WPIPE_Block2_start_1084_inst_req_0); -- 
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1084_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1084_Update/req
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1084_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1084_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1084_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1084_update_start_
      -- 
    ack_2355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1084_inst_ack_0, ack => convTranspose_CP_34_elements(303)); -- 
    req_2359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(303), ack => WPIPE_Block2_start_1084_inst_req_1); -- 
    -- CP-element group 304:  transition  input  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (6) 
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1084_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1087_Sample/$entry
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1084_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1087_sample_start_
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1084_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1087_Sample/req
      -- 
    ack_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1084_inst_ack_1, ack => convTranspose_CP_34_elements(304)); -- 
    req_2368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(304), ack => WPIPE_Block2_start_1087_inst_req_0); -- 
    -- CP-element group 305:  transition  input  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (6) 
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1087_update_start_
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1087_sample_completed_
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1087_Update/req
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1087_Update/$entry
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1087_Sample/ack
      -- CP-element group 305: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1087_Sample/$exit
      -- 
    ack_2369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1087_inst_ack_0, ack => convTranspose_CP_34_elements(305)); -- 
    req_2373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(305), ack => WPIPE_Block2_start_1087_inst_req_1); -- 
    -- CP-element group 306:  transition  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (6) 
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1087_update_completed_
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1090_Sample/req
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1087_Update/ack
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1090_Sample/$entry
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1087_Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1090_sample_start_
      -- 
    ack_2374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1087_inst_ack_1, ack => convTranspose_CP_34_elements(306)); -- 
    req_2382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(306), ack => WPIPE_Block2_start_1090_inst_req_0); -- 
    -- CP-element group 307:  transition  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1090_Update/req
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1090_Update/$entry
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1090_Sample/ack
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1090_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1090_update_start_
      -- CP-element group 307: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1090_sample_completed_
      -- 
    ack_2383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1090_inst_ack_0, ack => convTranspose_CP_34_elements(307)); -- 
    req_2387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(307), ack => WPIPE_Block2_start_1090_inst_req_1); -- 
    -- CP-element group 308:  transition  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (6) 
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1090_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1093_Sample/req
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1093_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1090_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1093_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1090_Update/ack
      -- 
    ack_2388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1090_inst_ack_1, ack => convTranspose_CP_34_elements(308)); -- 
    req_2396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(308), ack => WPIPE_Block2_start_1093_inst_req_0); -- 
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (6) 
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1093_Sample/$exit
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1093_update_start_
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1093_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1093_Sample/ack
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1093_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1093_Update/req
      -- 
    ack_2397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1093_inst_ack_0, ack => convTranspose_CP_34_elements(309)); -- 
    req_2401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(309), ack => WPIPE_Block2_start_1093_inst_req_1); -- 
    -- CP-element group 310:  transition  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (6) 
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1093_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1093_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1093_Update/ack
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1096_sample_start_
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1096_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1096_Sample/req
      -- 
    ack_2402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1093_inst_ack_1, ack => convTranspose_CP_34_elements(310)); -- 
    req_2410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(310), ack => WPIPE_Block2_start_1096_inst_req_0); -- 
    -- CP-element group 311:  transition  input  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (6) 
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1096_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1096_update_start_
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1096_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1096_Sample/ack
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1096_Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1096_Update/req
      -- 
    ack_2411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1096_inst_ack_0, ack => convTranspose_CP_34_elements(311)); -- 
    req_2415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(311), ack => WPIPE_Block2_start_1096_inst_req_1); -- 
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (6) 
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1096_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1096_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1096_Update/ack
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1099_sample_start_
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1099_Sample/$entry
      -- CP-element group 312: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1099_Sample/req
      -- 
    ack_2416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1096_inst_ack_1, ack => convTranspose_CP_34_elements(312)); -- 
    req_2424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(312), ack => WPIPE_Block2_start_1099_inst_req_0); -- 
    -- CP-element group 313:  transition  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (6) 
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1099_sample_completed_
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1099_update_start_
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1099_Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1099_Sample/ack
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1099_Update/$entry
      -- CP-element group 313: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1099_Update/req
      -- 
    ack_2425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1099_inst_ack_0, ack => convTranspose_CP_34_elements(313)); -- 
    req_2429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(313), ack => WPIPE_Block2_start_1099_inst_req_1); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	317 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1099_update_completed_
      -- CP-element group 314: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1099_Update/$exit
      -- CP-element group 314: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1099_Update/ack
      -- 
    ack_2430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1099_inst_ack_1, ack => convTranspose_CP_34_elements(314)); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	234 
    -- CP-element group 315: successors 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1110_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1110_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1110_Sample/ra
      -- 
    ra_2439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1110_inst_ack_0, ack => convTranspose_CP_34_elements(315)); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	234 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	317 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1110_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1110_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1110_Update/ca
      -- 
    ca_2444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1110_inst_ack_1, ack => convTranspose_CP_34_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	314 
    -- CP-element group 317: 	316 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1112_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1112_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1112_Sample/req
      -- 
    req_2452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(317), ack => WPIPE_Block2_start_1112_inst_req_0); -- 
    convTranspose_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(314) & convTranspose_CP_34_elements(316);
      gj_convTranspose_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  transition  input  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (6) 
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1112_sample_completed_
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1112_update_start_
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1112_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1112_Sample/ack
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1112_Update/$entry
      -- CP-element group 318: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1112_Update/req
      -- 
    ack_2453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1112_inst_ack_0, ack => convTranspose_CP_34_elements(318)); -- 
    req_2457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(318), ack => WPIPE_Block2_start_1112_inst_req_1); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	322 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1112_update_completed_
      -- CP-element group 319: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1112_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1112_Update/ack
      -- 
    ack_2458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1112_inst_ack_1, ack => convTranspose_CP_34_elements(319)); -- 
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	234 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1117_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1117_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1117_Sample/ra
      -- 
    ra_2467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1117_inst_ack_0, ack => convTranspose_CP_34_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	234 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1117_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1117_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1117_Update/ca
      -- 
    ca_2472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1117_inst_ack_1, ack => convTranspose_CP_34_elements(321)); -- 
    -- CP-element group 322:  join  transition  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	319 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1119_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1119_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1119_Sample/req
      -- 
    req_2480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(322), ack => WPIPE_Block2_start_1119_inst_req_0); -- 
    convTranspose_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(319) & convTranspose_CP_34_elements(321);
      gj_convTranspose_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  transition  input  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	322 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (6) 
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1119_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1119_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1119_update_start_
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1119_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1119_Sample/ack
      -- CP-element group 323: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1119_Update/req
      -- 
    ack_2481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1119_inst_ack_0, ack => convTranspose_CP_34_elements(323)); -- 
    req_2485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(323), ack => WPIPE_Block2_start_1119_inst_req_1); -- 
    -- CP-element group 324:  transition  input  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (6) 
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1119_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1119_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1119_Update/ack
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1122_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1122_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1122_Sample/req
      -- 
    ack_2486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1119_inst_ack_1, ack => convTranspose_CP_34_elements(324)); -- 
    req_2494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(324), ack => WPIPE_Block2_start_1122_inst_req_0); -- 
    -- CP-element group 325:  transition  input  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (6) 
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1122_sample_completed_
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1122_update_start_
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1122_Sample/$exit
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1122_Sample/ack
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1122_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1122_Update/req
      -- 
    ack_2495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1122_inst_ack_0, ack => convTranspose_CP_34_elements(325)); -- 
    req_2499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(325), ack => WPIPE_Block2_start_1122_inst_req_1); -- 
    -- CP-element group 326:  transition  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (6) 
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1122_update_completed_
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1122_Update/$exit
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1122_Update/ack
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1125_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1125_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1125_Sample/req
      -- 
    ack_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1122_inst_ack_1, ack => convTranspose_CP_34_elements(326)); -- 
    req_2508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(326), ack => WPIPE_Block2_start_1125_inst_req_0); -- 
    -- CP-element group 327:  transition  input  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (6) 
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1125_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1125_update_start_
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1125_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1125_Sample/ack
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1125_Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1125_Update/req
      -- 
    ack_2509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1125_inst_ack_0, ack => convTranspose_CP_34_elements(327)); -- 
    req_2513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(327), ack => WPIPE_Block2_start_1125_inst_req_1); -- 
    -- CP-element group 328:  transition  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (6) 
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1125_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1125_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1125_Update/ack
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1128_sample_start_
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1128_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1128_Sample/req
      -- 
    ack_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1125_inst_ack_1, ack => convTranspose_CP_34_elements(328)); -- 
    req_2522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(328), ack => WPIPE_Block2_start_1128_inst_req_0); -- 
    -- CP-element group 329:  transition  input  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329:  members (6) 
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1128_sample_completed_
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1128_update_start_
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1128_Sample/$exit
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1128_Sample/ack
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1128_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1128_Update/req
      -- 
    ack_2523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1128_inst_ack_0, ack => convTranspose_CP_34_elements(329)); -- 
    req_2527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(329), ack => WPIPE_Block2_start_1128_inst_req_1); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	373 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1128_update_completed_
      -- CP-element group 330: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1128_Update/$exit
      -- CP-element group 330: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block2_start_1128_Update/ack
      -- 
    ack_2528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1128_inst_ack_1, ack => convTranspose_CP_34_elements(330)); -- 
    -- CP-element group 331:  transition  input  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	234 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (6) 
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1131_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1131_update_start_
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1131_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1131_Sample/ack
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1131_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1131_Update/req
      -- 
    ack_2537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1131_inst_ack_0, ack => convTranspose_CP_34_elements(331)); -- 
    req_2541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(331), ack => WPIPE_Block3_start_1131_inst_req_1); -- 
    -- CP-element group 332:  transition  input  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (6) 
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1131_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1131_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1131_Update/ack
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1134_sample_start_
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1134_Sample/$entry
      -- CP-element group 332: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1134_Sample/req
      -- 
    ack_2542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1131_inst_ack_1, ack => convTranspose_CP_34_elements(332)); -- 
    req_2550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(332), ack => WPIPE_Block3_start_1134_inst_req_0); -- 
    -- CP-element group 333:  transition  input  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (6) 
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1134_sample_completed_
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1134_update_start_
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1134_Sample/$exit
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1134_Sample/ack
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1134_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1134_Update/req
      -- 
    ack_2551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1134_inst_ack_0, ack => convTranspose_CP_34_elements(333)); -- 
    req_2555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(333), ack => WPIPE_Block3_start_1134_inst_req_1); -- 
    -- CP-element group 334:  transition  input  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (6) 
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1134_update_completed_
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1134_Update/$exit
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1134_Update/ack
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1137_sample_start_
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1137_Sample/$entry
      -- CP-element group 334: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1137_Sample/req
      -- 
    ack_2556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1134_inst_ack_1, ack => convTranspose_CP_34_elements(334)); -- 
    req_2564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(334), ack => WPIPE_Block3_start_1137_inst_req_0); -- 
    -- CP-element group 335:  transition  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335:  members (6) 
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1137_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1137_update_start_
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1137_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1137_Sample/ack
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1137_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1137_Update/req
      -- 
    ack_2565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1137_inst_ack_0, ack => convTranspose_CP_34_elements(335)); -- 
    req_2569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(335), ack => WPIPE_Block3_start_1137_inst_req_1); -- 
    -- CP-element group 336:  transition  input  output  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	337 
    -- CP-element group 336:  members (6) 
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1137_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1137_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1137_Update/ack
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1140_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1140_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1140_Sample/req
      -- 
    ack_2570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1137_inst_ack_1, ack => convTranspose_CP_34_elements(336)); -- 
    req_2578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(336), ack => WPIPE_Block3_start_1140_inst_req_0); -- 
    -- CP-element group 337:  transition  input  output  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	336 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (6) 
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1140_sample_completed_
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1140_update_start_
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1140_Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1140_Sample/ack
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1140_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1140_Update/req
      -- 
    ack_2579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1140_inst_ack_0, ack => convTranspose_CP_34_elements(337)); -- 
    req_2583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(337), ack => WPIPE_Block3_start_1140_inst_req_1); -- 
    -- CP-element group 338:  transition  input  output  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (6) 
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1140_update_completed_
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1140_Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1140_Update/ack
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1143_sample_start_
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1143_Sample/$entry
      -- CP-element group 338: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1143_Sample/req
      -- 
    ack_2584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1140_inst_ack_1, ack => convTranspose_CP_34_elements(338)); -- 
    req_2592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(338), ack => WPIPE_Block3_start_1143_inst_req_0); -- 
    -- CP-element group 339:  transition  input  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (6) 
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1143_sample_completed_
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1143_update_start_
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1143_Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1143_Sample/ack
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1143_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1143_Update/req
      -- 
    ack_2593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1143_inst_ack_0, ack => convTranspose_CP_34_elements(339)); -- 
    req_2597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(339), ack => WPIPE_Block3_start_1143_inst_req_1); -- 
    -- CP-element group 340:  transition  input  output  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (6) 
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1143_update_completed_
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1143_Update/$exit
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1143_Update/ack
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1146_sample_start_
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1146_Sample/$entry
      -- CP-element group 340: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1146_Sample/req
      -- 
    ack_2598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1143_inst_ack_1, ack => convTranspose_CP_34_elements(340)); -- 
    req_2606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(340), ack => WPIPE_Block3_start_1146_inst_req_0); -- 
    -- CP-element group 341:  transition  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (6) 
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1146_sample_completed_
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1146_update_start_
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1146_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1146_Sample/ack
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1146_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1146_Update/req
      -- 
    ack_2607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1146_inst_ack_0, ack => convTranspose_CP_34_elements(341)); -- 
    req_2611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(341), ack => WPIPE_Block3_start_1146_inst_req_1); -- 
    -- CP-element group 342:  transition  input  output  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	343 
    -- CP-element group 342:  members (6) 
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1146_update_completed_
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1146_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1146_Update/ack
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1149_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1149_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1149_Sample/req
      -- 
    ack_2612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1146_inst_ack_1, ack => convTranspose_CP_34_elements(342)); -- 
    req_2620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(342), ack => WPIPE_Block3_start_1149_inst_req_0); -- 
    -- CP-element group 343:  transition  input  output  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	342 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (6) 
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1149_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1149_update_start_
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1149_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1149_Sample/ack
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1149_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1149_Update/req
      -- 
    ack_2621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1149_inst_ack_0, ack => convTranspose_CP_34_elements(343)); -- 
    req_2625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(343), ack => WPIPE_Block3_start_1149_inst_req_1); -- 
    -- CP-element group 344:  transition  input  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	345 
    -- CP-element group 344:  members (6) 
      -- CP-element group 344: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1149_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1149_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1149_Update/ack
      -- CP-element group 344: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1152_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1152_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1152_Sample/req
      -- 
    ack_2626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1149_inst_ack_1, ack => convTranspose_CP_34_elements(344)); -- 
    req_2634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(344), ack => WPIPE_Block3_start_1152_inst_req_0); -- 
    -- CP-element group 345:  transition  input  output  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	344 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345:  members (6) 
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1152_sample_completed_
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1152_update_start_
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1152_Sample/$exit
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1152_Sample/ack
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1152_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1152_Update/req
      -- 
    ack_2635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1152_inst_ack_0, ack => convTranspose_CP_34_elements(345)); -- 
    req_2639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(345), ack => WPIPE_Block3_start_1152_inst_req_1); -- 
    -- CP-element group 346:  transition  input  output  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (6) 
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1152_update_completed_
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1152_Update/$exit
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1152_Update/ack
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1155_sample_start_
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1155_Sample/$entry
      -- CP-element group 346: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1155_Sample/req
      -- 
    ack_2640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1152_inst_ack_1, ack => convTranspose_CP_34_elements(346)); -- 
    req_2648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(346), ack => WPIPE_Block3_start_1155_inst_req_0); -- 
    -- CP-element group 347:  transition  input  output  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (6) 
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1155_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1155_update_start_
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1155_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1155_Sample/ack
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1155_Update/$entry
      -- CP-element group 347: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1155_Update/req
      -- 
    ack_2649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1155_inst_ack_0, ack => convTranspose_CP_34_elements(347)); -- 
    req_2653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(347), ack => WPIPE_Block3_start_1155_inst_req_1); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	351 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1155_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1155_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1155_Update/ack
      -- 
    ack_2654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1155_inst_ack_1, ack => convTranspose_CP_34_elements(348)); -- 
    -- CP-element group 349:  transition  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	234 
    -- CP-element group 349: successors 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1166_sample_completed_
      -- CP-element group 349: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1166_Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1166_Sample/ra
      -- 
    ra_2663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1166_inst_ack_0, ack => convTranspose_CP_34_elements(349)); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	234 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1166_update_completed_
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1166_Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1166_Update/ca
      -- 
    ca_2668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1166_inst_ack_1, ack => convTranspose_CP_34_elements(350)); -- 
    -- CP-element group 351:  join  transition  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	348 
    -- CP-element group 351: 	350 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1168_sample_start_
      -- CP-element group 351: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1168_Sample/$entry
      -- CP-element group 351: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1168_Sample/req
      -- 
    req_2676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(351), ack => WPIPE_Block3_start_1168_inst_req_0); -- 
    convTranspose_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(348) & convTranspose_CP_34_elements(350);
      gj_convTranspose_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  transition  input  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (6) 
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1168_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1168_update_start_
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1168_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1168_Sample/ack
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1168_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1168_Update/req
      -- 
    ack_2677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1168_inst_ack_0, ack => convTranspose_CP_34_elements(352)); -- 
    req_2681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(352), ack => WPIPE_Block3_start_1168_inst_req_1); -- 
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	356 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1168_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1168_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1168_Update/ack
      -- 
    ack_2682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1168_inst_ack_1, ack => convTranspose_CP_34_elements(353)); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	234 
    -- CP-element group 354: successors 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1173_sample_completed_
      -- CP-element group 354: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1173_Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1173_Sample/ra
      -- 
    ra_2691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1173_inst_ack_0, ack => convTranspose_CP_34_elements(354)); -- 
    -- CP-element group 355:  transition  input  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	234 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1173_update_completed_
      -- CP-element group 355: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1173_Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/type_cast_1173_Update/ca
      -- 
    ca_2696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1173_inst_ack_1, ack => convTranspose_CP_34_elements(355)); -- 
    -- CP-element group 356:  join  transition  output  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	353 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1175_sample_start_
      -- CP-element group 356: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1175_Sample/$entry
      -- CP-element group 356: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1175_Sample/req
      -- 
    req_2704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(356), ack => WPIPE_Block3_start_1175_inst_req_0); -- 
    convTranspose_cp_element_group_356: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_356"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(353) & convTranspose_CP_34_elements(355);
      gj_convTranspose_cp_element_group_356 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(356), clk => clk, reset => reset); --
    end block;
    -- CP-element group 357:  transition  input  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (6) 
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1175_sample_completed_
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1175_update_start_
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1175_Sample/$exit
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1175_Sample/ack
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1175_Update/$entry
      -- CP-element group 357: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1175_Update/req
      -- 
    ack_2705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1175_inst_ack_0, ack => convTranspose_CP_34_elements(357)); -- 
    req_2709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(357), ack => WPIPE_Block3_start_1175_inst_req_1); -- 
    -- CP-element group 358:  transition  input  output  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (6) 
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1175_update_completed_
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1175_Update/$exit
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1175_Update/ack
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1178_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1178_Sample/$entry
      -- CP-element group 358: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1178_Sample/req
      -- 
    ack_2710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1175_inst_ack_1, ack => convTranspose_CP_34_elements(358)); -- 
    req_2718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(358), ack => WPIPE_Block3_start_1178_inst_req_0); -- 
    -- CP-element group 359:  transition  input  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (6) 
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1178_sample_completed_
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1178_update_start_
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1178_Sample/$exit
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1178_Sample/ack
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1178_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1178_Update/req
      -- 
    ack_2719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1178_inst_ack_0, ack => convTranspose_CP_34_elements(359)); -- 
    req_2723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(359), ack => WPIPE_Block3_start_1178_inst_req_1); -- 
    -- CP-element group 360:  transition  input  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360:  members (6) 
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1178_update_completed_
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1178_Update/$exit
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1178_Update/ack
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1181_sample_start_
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1181_Sample/$entry
      -- CP-element group 360: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1181_Sample/req
      -- 
    ack_2724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1178_inst_ack_1, ack => convTranspose_CP_34_elements(360)); -- 
    req_2732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(360), ack => WPIPE_Block3_start_1181_inst_req_0); -- 
    -- CP-element group 361:  transition  input  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (6) 
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1181_sample_completed_
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1181_update_start_
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1181_Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1181_Sample/ack
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1181_Update/$entry
      -- CP-element group 361: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1181_Update/req
      -- 
    ack_2733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1181_inst_ack_0, ack => convTranspose_CP_34_elements(361)); -- 
    req_2737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(361), ack => WPIPE_Block3_start_1181_inst_req_1); -- 
    -- CP-element group 362:  transition  input  output  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (6) 
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1181_update_completed_
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1181_Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1181_Update/ack
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1184_sample_start_
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1184_Sample/$entry
      -- CP-element group 362: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1184_Sample/req
      -- 
    ack_2738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1181_inst_ack_1, ack => convTranspose_CP_34_elements(362)); -- 
    req_2746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(362), ack => WPIPE_Block3_start_1184_inst_req_0); -- 
    -- CP-element group 363:  transition  input  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (6) 
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1184_sample_completed_
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1184_update_start_
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1184_Sample/$exit
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1184_Sample/ack
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1184_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1184_Update/req
      -- 
    ack_2747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1184_inst_ack_0, ack => convTranspose_CP_34_elements(363)); -- 
    req_2751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(363), ack => WPIPE_Block3_start_1184_inst_req_1); -- 
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	373 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1184_update_completed_
      -- CP-element group 364: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1184_Update/$exit
      -- CP-element group 364: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/WPIPE_Block3_start_1184_Update/ack
      -- 
    ack_2752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1184_inst_ack_1, ack => convTranspose_CP_34_elements(364)); -- 
    -- CP-element group 365:  transition  input  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	234 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (6) 
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block0_done_1188_sample_completed_
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block0_done_1188_update_start_
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block0_done_1188_Sample/$exit
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block0_done_1188_Sample/ra
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block0_done_1188_Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block0_done_1188_Update/cr
      -- 
    ra_2761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1188_inst_ack_0, ack => convTranspose_CP_34_elements(365)); -- 
    cr_2765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(365), ack => RPIPE_Block0_done_1188_inst_req_1); -- 
    -- CP-element group 366:  transition  input  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	373 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block0_done_1188_update_completed_
      -- CP-element group 366: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block0_done_1188_Update/$exit
      -- CP-element group 366: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block0_done_1188_Update/ca
      -- 
    ca_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1188_inst_ack_1, ack => convTranspose_CP_34_elements(366)); -- 
    -- CP-element group 367:  transition  input  output  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	234 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (6) 
      -- CP-element group 367: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block1_done_1191_sample_completed_
      -- CP-element group 367: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block1_done_1191_update_start_
      -- CP-element group 367: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block1_done_1191_Sample/$exit
      -- CP-element group 367: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block1_done_1191_Sample/ra
      -- CP-element group 367: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block1_done_1191_Update/$entry
      -- CP-element group 367: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block1_done_1191_Update/cr
      -- 
    ra_2775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1191_inst_ack_0, ack => convTranspose_CP_34_elements(367)); -- 
    cr_2779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(367), ack => RPIPE_Block1_done_1191_inst_req_1); -- 
    -- CP-element group 368:  transition  input  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	373 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block1_done_1191_update_completed_
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block1_done_1191_Update/$exit
      -- CP-element group 368: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block1_done_1191_Update/ca
      -- 
    ca_2780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1191_inst_ack_1, ack => convTranspose_CP_34_elements(368)); -- 
    -- CP-element group 369:  transition  input  output  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	234 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (6) 
      -- CP-element group 369: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block2_done_1194_sample_completed_
      -- CP-element group 369: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block2_done_1194_update_start_
      -- CP-element group 369: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block2_done_1194_Sample/$exit
      -- CP-element group 369: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block2_done_1194_Sample/ra
      -- CP-element group 369: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block2_done_1194_Update/$entry
      -- CP-element group 369: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block2_done_1194_Update/cr
      -- 
    ra_2789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1194_inst_ack_0, ack => convTranspose_CP_34_elements(369)); -- 
    cr_2793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(369), ack => RPIPE_Block2_done_1194_inst_req_1); -- 
    -- CP-element group 370:  transition  input  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	373 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block2_done_1194_update_completed_
      -- CP-element group 370: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block2_done_1194_Update/$exit
      -- CP-element group 370: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block2_done_1194_Update/ca
      -- 
    ca_2794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1194_inst_ack_1, ack => convTranspose_CP_34_elements(370)); -- 
    -- CP-element group 371:  transition  input  output  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	234 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (6) 
      -- CP-element group 371: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block3_done_1197_sample_completed_
      -- CP-element group 371: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block3_done_1197_update_start_
      -- CP-element group 371: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block3_done_1197_Sample/$exit
      -- CP-element group 371: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block3_done_1197_Sample/ra
      -- CP-element group 371: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block3_done_1197_Update/$entry
      -- CP-element group 371: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block3_done_1197_Update/cr
      -- 
    ra_2803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1197_inst_ack_0, ack => convTranspose_CP_34_elements(371)); -- 
    cr_2807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(371), ack => RPIPE_Block3_done_1197_inst_req_1); -- 
    -- CP-element group 372:  transition  input  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block3_done_1197_update_completed_
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block3_done_1197_Update/$exit
      -- CP-element group 372: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/RPIPE_Block3_done_1197_Update/ca
      -- 
    ca_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1197_inst_ack_1, ack => convTranspose_CP_34_elements(372)); -- 
    -- CP-element group 373:  join  fork  transition  place  output  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	262 
    -- CP-element group 373: 	296 
    -- CP-element group 373: 	330 
    -- CP-element group 373: 	364 
    -- CP-element group 373: 	366 
    -- CP-element group 373: 	368 
    -- CP-element group 373: 	370 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373: 	375 
    -- CP-element group 373: 	377 
    -- CP-element group 373: 	379 
    -- CP-element group 373: 	381 
    -- CP-element group 373: 	383 
    -- CP-element group 373: 	385 
    -- CP-element group 373: 	387 
    -- CP-element group 373: 	389 
    -- CP-element group 373: 	391 
    -- CP-element group 373: 	393 
    -- CP-element group 373:  members (37) 
      -- CP-element group 373: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198__exit__
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309__entry__
      -- CP-element group 373: 	 branch_block_stmt_38/assign_stmt_977_to_assign_stmt_1198/$exit
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/$entry
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/call_stmt_1201_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/call_stmt_1201_update_start_
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/call_stmt_1201_Sample/$entry
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/call_stmt_1201_Sample/crr
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/call_stmt_1201_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/call_stmt_1201_Update/ccr
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1205_update_start_
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1205_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1205_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1214_update_start_
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1214_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1214_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1224_update_start_
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1224_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1224_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1234_update_start_
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1234_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1234_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1244_update_start_
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1244_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1244_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1254_update_start_
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1254_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1254_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1264_update_start_
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1264_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1264_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1274_update_start_
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1274_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1274_Update/cr
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1284_update_start_
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1284_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1284_Update/cr
      -- 
    crr_2819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(373), ack => call_stmt_1201_call_req_0); -- 
    ccr_2824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(373), ack => call_stmt_1201_call_req_1); -- 
    cr_2838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(373), ack => type_cast_1205_inst_req_1); -- 
    cr_2852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(373), ack => type_cast_1214_inst_req_1); -- 
    cr_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(373), ack => type_cast_1224_inst_req_1); -- 
    cr_2880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(373), ack => type_cast_1234_inst_req_1); -- 
    cr_2894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(373), ack => type_cast_1244_inst_req_1); -- 
    cr_2908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(373), ack => type_cast_1254_inst_req_1); -- 
    cr_2922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(373), ack => type_cast_1264_inst_req_1); -- 
    cr_2936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(373), ack => type_cast_1274_inst_req_1); -- 
    cr_2950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(373), ack => type_cast_1284_inst_req_1); -- 
    convTranspose_cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_373"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(262) & convTranspose_CP_34_elements(296) & convTranspose_CP_34_elements(330) & convTranspose_CP_34_elements(364) & convTranspose_CP_34_elements(366) & convTranspose_CP_34_elements(368) & convTranspose_CP_34_elements(370) & convTranspose_CP_34_elements(372);
      gj_convTranspose_cp_element_group_373 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 374:  transition  input  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/call_stmt_1201_sample_completed_
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/call_stmt_1201_Sample/$exit
      -- CP-element group 374: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/call_stmt_1201_Sample/cra
      -- 
    cra_2820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1201_call_ack_0, ack => convTranspose_CP_34_elements(374)); -- 
    -- CP-element group 375:  transition  input  output  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	373 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375:  members (6) 
      -- CP-element group 375: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/call_stmt_1201_update_completed_
      -- CP-element group 375: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/call_stmt_1201_Update/$exit
      -- CP-element group 375: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/call_stmt_1201_Update/cca
      -- CP-element group 375: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1205_sample_start_
      -- CP-element group 375: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1205_Sample/$entry
      -- CP-element group 375: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1205_Sample/rr
      -- 
    cca_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1201_call_ack_1, ack => convTranspose_CP_34_elements(375)); -- 
    rr_2833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(375), ack => type_cast_1205_inst_req_0); -- 
    -- CP-element group 376:  transition  input  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	375 
    -- CP-element group 376: successors 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1205_sample_completed_
      -- CP-element group 376: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1205_Sample/$exit
      -- CP-element group 376: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1205_Sample/ra
      -- 
    ra_2834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1205_inst_ack_0, ack => convTranspose_CP_34_elements(376)); -- 
    -- CP-element group 377:  fork  transition  input  output  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	373 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	378 
    -- CP-element group 377: 	380 
    -- CP-element group 377: 	382 
    -- CP-element group 377: 	384 
    -- CP-element group 377: 	386 
    -- CP-element group 377: 	388 
    -- CP-element group 377: 	390 
    -- CP-element group 377: 	392 
    -- CP-element group 377:  members (27) 
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1205_update_completed_
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1205_Update/$exit
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1205_Update/ca
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1214_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1214_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1214_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1224_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1224_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1224_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1234_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1234_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1234_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1244_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1244_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1244_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1254_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1254_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1254_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1264_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1264_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1264_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1274_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1274_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1274_Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1284_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1284_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1284_Sample/rr
      -- 
    ca_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1205_inst_ack_1, ack => convTranspose_CP_34_elements(377)); -- 
    rr_2847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(377), ack => type_cast_1214_inst_req_0); -- 
    rr_2861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(377), ack => type_cast_1224_inst_req_0); -- 
    rr_2875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(377), ack => type_cast_1234_inst_req_0); -- 
    rr_2889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(377), ack => type_cast_1244_inst_req_0); -- 
    rr_2903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(377), ack => type_cast_1254_inst_req_0); -- 
    rr_2917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(377), ack => type_cast_1264_inst_req_0); -- 
    rr_2931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(377), ack => type_cast_1274_inst_req_0); -- 
    rr_2945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(377), ack => type_cast_1284_inst_req_0); -- 
    -- CP-element group 378:  transition  input  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	377 
    -- CP-element group 378: successors 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1214_sample_completed_
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1214_Sample/$exit
      -- CP-element group 378: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1214_Sample/ra
      -- 
    ra_2848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1214_inst_ack_0, ack => convTranspose_CP_34_elements(378)); -- 
    -- CP-element group 379:  transition  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	373 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	414 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1214_update_completed_
      -- CP-element group 379: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1214_Update/$exit
      -- CP-element group 379: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1214_Update/ca
      -- 
    ca_2853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1214_inst_ack_1, ack => convTranspose_CP_34_elements(379)); -- 
    -- CP-element group 380:  transition  input  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	377 
    -- CP-element group 380: successors 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1224_sample_completed_
      -- CP-element group 380: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1224_Sample/$exit
      -- CP-element group 380: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1224_Sample/ra
      -- 
    ra_2862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1224_inst_ack_0, ack => convTranspose_CP_34_elements(380)); -- 
    -- CP-element group 381:  transition  input  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	373 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	411 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1224_update_completed_
      -- CP-element group 381: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1224_Update/$exit
      -- CP-element group 381: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1224_Update/ca
      -- 
    ca_2867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1224_inst_ack_1, ack => convTranspose_CP_34_elements(381)); -- 
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	377 
    -- CP-element group 382: successors 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1234_sample_completed_
      -- CP-element group 382: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1234_Sample/$exit
      -- CP-element group 382: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1234_Sample/ra
      -- 
    ra_2876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1234_inst_ack_0, ack => convTranspose_CP_34_elements(382)); -- 
    -- CP-element group 383:  transition  input  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	373 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	408 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1234_update_completed_
      -- CP-element group 383: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1234_Update/$exit
      -- CP-element group 383: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1234_Update/ca
      -- 
    ca_2881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1234_inst_ack_1, ack => convTranspose_CP_34_elements(383)); -- 
    -- CP-element group 384:  transition  input  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	377 
    -- CP-element group 384: successors 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1244_sample_completed_
      -- CP-element group 384: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1244_Sample/$exit
      -- CP-element group 384: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1244_Sample/ra
      -- 
    ra_2890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1244_inst_ack_0, ack => convTranspose_CP_34_elements(384)); -- 
    -- CP-element group 385:  transition  input  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	373 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	405 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1244_update_completed_
      -- CP-element group 385: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1244_Update/$exit
      -- CP-element group 385: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1244_Update/ca
      -- 
    ca_2895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1244_inst_ack_1, ack => convTranspose_CP_34_elements(385)); -- 
    -- CP-element group 386:  transition  input  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	377 
    -- CP-element group 386: successors 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1254_sample_completed_
      -- CP-element group 386: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1254_Sample/$exit
      -- CP-element group 386: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1254_Sample/ra
      -- 
    ra_2904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1254_inst_ack_0, ack => convTranspose_CP_34_elements(386)); -- 
    -- CP-element group 387:  transition  input  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	373 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	402 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1254_update_completed_
      -- CP-element group 387: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1254_Update/$exit
      -- CP-element group 387: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1254_Update/ca
      -- 
    ca_2909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1254_inst_ack_1, ack => convTranspose_CP_34_elements(387)); -- 
    -- CP-element group 388:  transition  input  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	377 
    -- CP-element group 388: successors 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1264_sample_completed_
      -- CP-element group 388: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1264_Sample/$exit
      -- CP-element group 388: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1264_Sample/ra
      -- 
    ra_2918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1264_inst_ack_0, ack => convTranspose_CP_34_elements(388)); -- 
    -- CP-element group 389:  transition  input  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	373 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	399 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1264_update_completed_
      -- CP-element group 389: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1264_Update/$exit
      -- CP-element group 389: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1264_Update/ca
      -- 
    ca_2923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1264_inst_ack_1, ack => convTranspose_CP_34_elements(389)); -- 
    -- CP-element group 390:  transition  input  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	377 
    -- CP-element group 390: successors 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1274_sample_completed_
      -- CP-element group 390: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1274_Sample/$exit
      -- CP-element group 390: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1274_Sample/ra
      -- 
    ra_2932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1274_inst_ack_0, ack => convTranspose_CP_34_elements(390)); -- 
    -- CP-element group 391:  transition  input  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	373 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	396 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1274_update_completed_
      -- CP-element group 391: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1274_Update/$exit
      -- CP-element group 391: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1274_Update/ca
      -- 
    ca_2937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1274_inst_ack_1, ack => convTranspose_CP_34_elements(391)); -- 
    -- CP-element group 392:  transition  input  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	377 
    -- CP-element group 392: successors 
    -- CP-element group 392:  members (3) 
      -- CP-element group 392: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1284_sample_completed_
      -- CP-element group 392: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1284_Sample/$exit
      -- CP-element group 392: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1284_Sample/ra
      -- 
    ra_2946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1284_inst_ack_0, ack => convTranspose_CP_34_elements(392)); -- 
    -- CP-element group 393:  transition  input  output  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	373 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	394 
    -- CP-element group 393:  members (6) 
      -- CP-element group 393: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1284_update_completed_
      -- CP-element group 393: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1284_Update/$exit
      -- CP-element group 393: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/type_cast_1284_Update/ca
      -- CP-element group 393: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1286_sample_start_
      -- CP-element group 393: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1286_Sample/$entry
      -- CP-element group 393: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1286_Sample/req
      -- 
    ca_2951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1284_inst_ack_1, ack => convTranspose_CP_34_elements(393)); -- 
    req_2959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(393), ack => WPIPE_ConvTranspose_output_pipe_1286_inst_req_0); -- 
    -- CP-element group 394:  transition  input  output  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	393 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	395 
    -- CP-element group 394:  members (6) 
      -- CP-element group 394: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1286_Update/req
      -- CP-element group 394: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1286_Update/$entry
      -- CP-element group 394: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1286_sample_completed_
      -- CP-element group 394: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1286_update_start_
      -- CP-element group 394: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1286_Sample/$exit
      -- CP-element group 394: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1286_Sample/ack
      -- 
    ack_2960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1286_inst_ack_0, ack => convTranspose_CP_34_elements(394)); -- 
    req_2964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(394), ack => WPIPE_ConvTranspose_output_pipe_1286_inst_req_1); -- 
    -- CP-element group 395:  transition  input  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	394 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	396 
    -- CP-element group 395:  members (3) 
      -- CP-element group 395: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1286_Update/ack
      -- CP-element group 395: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1286_Update/$exit
      -- CP-element group 395: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1286_update_completed_
      -- 
    ack_2965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1286_inst_ack_1, ack => convTranspose_CP_34_elements(395)); -- 
    -- CP-element group 396:  join  transition  output  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	391 
    -- CP-element group 396: 	395 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	397 
    -- CP-element group 396:  members (3) 
      -- CP-element group 396: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1289_sample_start_
      -- CP-element group 396: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1289_Sample/req
      -- CP-element group 396: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1289_Sample/$entry
      -- 
    req_2973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(396), ack => WPIPE_ConvTranspose_output_pipe_1289_inst_req_0); -- 
    convTranspose_cp_element_group_396: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_396"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(391) & convTranspose_CP_34_elements(395);
      gj_convTranspose_cp_element_group_396 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(396), clk => clk, reset => reset); --
    end block;
    -- CP-element group 397:  transition  input  output  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	396 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	398 
    -- CP-element group 397:  members (6) 
      -- CP-element group 397: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1289_sample_completed_
      -- CP-element group 397: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1289_Sample/$exit
      -- CP-element group 397: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1289_update_start_
      -- CP-element group 397: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1289_Sample/ack
      -- CP-element group 397: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1289_Update/$entry
      -- CP-element group 397: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1289_Update/req
      -- 
    ack_2974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1289_inst_ack_0, ack => convTranspose_CP_34_elements(397)); -- 
    req_2978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(397), ack => WPIPE_ConvTranspose_output_pipe_1289_inst_req_1); -- 
    -- CP-element group 398:  transition  input  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	397 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	399 
    -- CP-element group 398:  members (3) 
      -- CP-element group 398: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1289_Update/$exit
      -- CP-element group 398: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1289_update_completed_
      -- CP-element group 398: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1289_Update/ack
      -- 
    ack_2979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1289_inst_ack_1, ack => convTranspose_CP_34_elements(398)); -- 
    -- CP-element group 399:  join  transition  output  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	389 
    -- CP-element group 399: 	398 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	400 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1292_Sample/req
      -- CP-element group 399: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1292_Sample/$entry
      -- CP-element group 399: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1292_sample_start_
      -- 
    req_2987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(399), ack => WPIPE_ConvTranspose_output_pipe_1292_inst_req_0); -- 
    convTranspose_cp_element_group_399: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_399"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(389) & convTranspose_CP_34_elements(398);
      gj_convTranspose_cp_element_group_399 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(399), clk => clk, reset => reset); --
    end block;
    -- CP-element group 400:  transition  input  output  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	399 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	401 
    -- CP-element group 400:  members (6) 
      -- CP-element group 400: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1292_Update/req
      -- CP-element group 400: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1292_Update/$entry
      -- CP-element group 400: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1292_Sample/ack
      -- CP-element group 400: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1292_Sample/$exit
      -- CP-element group 400: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1292_update_start_
      -- CP-element group 400: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1292_sample_completed_
      -- 
    ack_2988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1292_inst_ack_0, ack => convTranspose_CP_34_elements(400)); -- 
    req_2992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(400), ack => WPIPE_ConvTranspose_output_pipe_1292_inst_req_1); -- 
    -- CP-element group 401:  transition  input  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	400 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	402 
    -- CP-element group 401:  members (3) 
      -- CP-element group 401: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1292_Update/ack
      -- CP-element group 401: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1292_Update/$exit
      -- CP-element group 401: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1292_update_completed_
      -- 
    ack_2993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1292_inst_ack_1, ack => convTranspose_CP_34_elements(401)); -- 
    -- CP-element group 402:  join  transition  output  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	387 
    -- CP-element group 402: 	401 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	403 
    -- CP-element group 402:  members (3) 
      -- CP-element group 402: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1295_Sample/req
      -- CP-element group 402: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1295_Sample/$entry
      -- CP-element group 402: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1295_sample_start_
      -- 
    req_3001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(402), ack => WPIPE_ConvTranspose_output_pipe_1295_inst_req_0); -- 
    convTranspose_cp_element_group_402: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_402"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(387) & convTranspose_CP_34_elements(401);
      gj_convTranspose_cp_element_group_402 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(402), clk => clk, reset => reset); --
    end block;
    -- CP-element group 403:  transition  input  output  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	402 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	404 
    -- CP-element group 403:  members (6) 
      -- CP-element group 403: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1295_Update/req
      -- CP-element group 403: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1295_Update/$entry
      -- CP-element group 403: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1295_Sample/ack
      -- CP-element group 403: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1295_Sample/$exit
      -- CP-element group 403: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1295_update_start_
      -- CP-element group 403: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1295_sample_completed_
      -- 
    ack_3002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1295_inst_ack_0, ack => convTranspose_CP_34_elements(403)); -- 
    req_3006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(403), ack => WPIPE_ConvTranspose_output_pipe_1295_inst_req_1); -- 
    -- CP-element group 404:  transition  input  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	403 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	405 
    -- CP-element group 404:  members (3) 
      -- CP-element group 404: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1295_Update/ack
      -- CP-element group 404: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1295_Update/$exit
      -- CP-element group 404: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1295_update_completed_
      -- 
    ack_3007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1295_inst_ack_1, ack => convTranspose_CP_34_elements(404)); -- 
    -- CP-element group 405:  join  transition  output  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	385 
    -- CP-element group 405: 	404 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	406 
    -- CP-element group 405:  members (3) 
      -- CP-element group 405: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1298_Sample/req
      -- CP-element group 405: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1298_Sample/$entry
      -- CP-element group 405: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1298_sample_start_
      -- 
    req_3015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(405), ack => WPIPE_ConvTranspose_output_pipe_1298_inst_req_0); -- 
    convTranspose_cp_element_group_405: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_405"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(385) & convTranspose_CP_34_elements(404);
      gj_convTranspose_cp_element_group_405 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(405), clk => clk, reset => reset); --
    end block;
    -- CP-element group 406:  transition  input  output  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	405 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	407 
    -- CP-element group 406:  members (6) 
      -- CP-element group 406: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1298_Sample/ack
      -- CP-element group 406: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1298_Update/req
      -- CP-element group 406: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1298_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1298_Sample/$exit
      -- CP-element group 406: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1298_update_start_
      -- CP-element group 406: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1298_sample_completed_
      -- 
    ack_3016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1298_inst_ack_0, ack => convTranspose_CP_34_elements(406)); -- 
    req_3020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(406), ack => WPIPE_ConvTranspose_output_pipe_1298_inst_req_1); -- 
    -- CP-element group 407:  transition  input  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	406 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	408 
    -- CP-element group 407:  members (3) 
      -- CP-element group 407: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1298_Update/ack
      -- CP-element group 407: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1298_Update/$exit
      -- CP-element group 407: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1298_update_completed_
      -- 
    ack_3021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1298_inst_ack_1, ack => convTranspose_CP_34_elements(407)); -- 
    -- CP-element group 408:  join  transition  output  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	383 
    -- CP-element group 408: 	407 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	409 
    -- CP-element group 408:  members (3) 
      -- CP-element group 408: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1301_Sample/$entry
      -- CP-element group 408: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1301_Sample/req
      -- CP-element group 408: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1301_sample_start_
      -- 
    req_3029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(408), ack => WPIPE_ConvTranspose_output_pipe_1301_inst_req_0); -- 
    convTranspose_cp_element_group_408: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_408"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(383) & convTranspose_CP_34_elements(407);
      gj_convTranspose_cp_element_group_408 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(408), clk => clk, reset => reset); --
    end block;
    -- CP-element group 409:  transition  input  output  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	408 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	410 
    -- CP-element group 409:  members (6) 
      -- CP-element group 409: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1301_Sample/ack
      -- CP-element group 409: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1301_Update/$entry
      -- CP-element group 409: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1301_Sample/$exit
      -- CP-element group 409: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1301_sample_completed_
      -- CP-element group 409: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1301_Update/req
      -- CP-element group 409: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1301_update_start_
      -- 
    ack_3030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1301_inst_ack_0, ack => convTranspose_CP_34_elements(409)); -- 
    req_3034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(409), ack => WPIPE_ConvTranspose_output_pipe_1301_inst_req_1); -- 
    -- CP-element group 410:  transition  input  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	409 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	411 
    -- CP-element group 410:  members (3) 
      -- CP-element group 410: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1301_Update/$exit
      -- CP-element group 410: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1301_Update/ack
      -- CP-element group 410: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1301_update_completed_
      -- 
    ack_3035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1301_inst_ack_1, ack => convTranspose_CP_34_elements(410)); -- 
    -- CP-element group 411:  join  transition  output  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	381 
    -- CP-element group 411: 	410 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	412 
    -- CP-element group 411:  members (3) 
      -- CP-element group 411: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1304_sample_start_
      -- CP-element group 411: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1304_Sample/req
      -- CP-element group 411: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1304_Sample/$entry
      -- 
    req_3043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(411), ack => WPIPE_ConvTranspose_output_pipe_1304_inst_req_0); -- 
    convTranspose_cp_element_group_411: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_411"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(381) & convTranspose_CP_34_elements(410);
      gj_convTranspose_cp_element_group_411 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(411), clk => clk, reset => reset); --
    end block;
    -- CP-element group 412:  transition  input  output  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	411 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	413 
    -- CP-element group 412:  members (6) 
      -- CP-element group 412: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1304_sample_completed_
      -- CP-element group 412: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1304_update_start_
      -- CP-element group 412: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1304_Update/req
      -- CP-element group 412: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1304_Update/$entry
      -- CP-element group 412: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1304_Sample/ack
      -- CP-element group 412: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1304_Sample/$exit
      -- 
    ack_3044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1304_inst_ack_0, ack => convTranspose_CP_34_elements(412)); -- 
    req_3048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(412), ack => WPIPE_ConvTranspose_output_pipe_1304_inst_req_1); -- 
    -- CP-element group 413:  transition  input  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	412 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	414 
    -- CP-element group 413:  members (3) 
      -- CP-element group 413: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1304_update_completed_
      -- CP-element group 413: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1304_Update/ack
      -- CP-element group 413: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1304_Update/$exit
      -- 
    ack_3049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1304_inst_ack_1, ack => convTranspose_CP_34_elements(413)); -- 
    -- CP-element group 414:  join  transition  output  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	379 
    -- CP-element group 414: 	413 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1307_Sample/req
      -- CP-element group 414: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1307_Sample/$entry
      -- CP-element group 414: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1307_sample_start_
      -- 
    req_3057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(414), ack => WPIPE_ConvTranspose_output_pipe_1307_inst_req_0); -- 
    convTranspose_cp_element_group_414: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_414"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(379) & convTranspose_CP_34_elements(413);
      gj_convTranspose_cp_element_group_414 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(414), clk => clk, reset => reset); --
    end block;
    -- CP-element group 415:  transition  input  output  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	414 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	416 
    -- CP-element group 415:  members (6) 
      -- CP-element group 415: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1307_Update/req
      -- CP-element group 415: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1307_Update/$entry
      -- CP-element group 415: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1307_Sample/ack
      -- CP-element group 415: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1307_Sample/$exit
      -- CP-element group 415: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1307_update_start_
      -- CP-element group 415: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1307_sample_completed_
      -- 
    ack_3058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 415_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1307_inst_ack_0, ack => convTranspose_CP_34_elements(415)); -- 
    req_3062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(415), ack => WPIPE_ConvTranspose_output_pipe_1307_inst_req_1); -- 
    -- CP-element group 416:  branch  transition  place  input  output  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	415 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	417 
    -- CP-element group 416: 	418 
    -- CP-element group 416:  members (13) 
      -- CP-element group 416: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309__exit__
      -- CP-element group 416: 	 branch_block_stmt_38/if_stmt_1311__entry__
      -- CP-element group 416: 	 branch_block_stmt_38/if_stmt_1311_else_link/$entry
      -- CP-element group 416: 	 branch_block_stmt_38/if_stmt_1311_if_link/$entry
      -- CP-element group 416: 	 branch_block_stmt_38/if_stmt_1311_eval_test/branch_req
      -- CP-element group 416: 	 branch_block_stmt_38/if_stmt_1311_eval_test/$exit
      -- CP-element group 416: 	 branch_block_stmt_38/if_stmt_1311_eval_test/$entry
      -- CP-element group 416: 	 branch_block_stmt_38/if_stmt_1311_dead_link/$entry
      -- CP-element group 416: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1307_Update/ack
      -- CP-element group 416: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1307_Update/$exit
      -- CP-element group 416: 	 branch_block_stmt_38/R_cmp264505_1312_place
      -- CP-element group 416: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/WPIPE_ConvTranspose_output_pipe_1307_update_completed_
      -- CP-element group 416: 	 branch_block_stmt_38/call_stmt_1201_to_assign_stmt_1309/$exit
      -- 
    ack_3063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1307_inst_ack_1, ack => convTranspose_CP_34_elements(416)); -- 
    branch_req_3071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(416), ack => if_stmt_1311_branch_req_0); -- 
    -- CP-element group 417:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	416 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	419 
    -- CP-element group 417: 	420 
    -- CP-element group 417:  members (18) 
      -- CP-element group 417: 	 branch_block_stmt_38/merge_stmt_1317__exit__
      -- CP-element group 417: 	 branch_block_stmt_38/assign_stmt_1323_to_assign_stmt_1352__entry__
      -- CP-element group 417: 	 branch_block_stmt_38/assign_stmt_1323_to_assign_stmt_1352/type_cast_1338_Update/cr
      -- CP-element group 417: 	 branch_block_stmt_38/assign_stmt_1323_to_assign_stmt_1352/type_cast_1338_Update/$entry
      -- CP-element group 417: 	 branch_block_stmt_38/assign_stmt_1323_to_assign_stmt_1352/type_cast_1338_Sample/rr
      -- CP-element group 417: 	 branch_block_stmt_38/assign_stmt_1323_to_assign_stmt_1352/type_cast_1338_Sample/$entry
      -- CP-element group 417: 	 branch_block_stmt_38/assign_stmt_1323_to_assign_stmt_1352/type_cast_1338_update_start_
      -- CP-element group 417: 	 branch_block_stmt_38/assign_stmt_1323_to_assign_stmt_1352/type_cast_1338_sample_start_
      -- CP-element group 417: 	 branch_block_stmt_38/assign_stmt_1323_to_assign_stmt_1352/$entry
      -- CP-element group 417: 	 branch_block_stmt_38/if_stmt_1311_if_link/if_choice_transition
      -- CP-element group 417: 	 branch_block_stmt_38/if_stmt_1311_if_link/$exit
      -- CP-element group 417: 	 branch_block_stmt_38/forx_xend273_bbx_xnph
      -- CP-element group 417: 	 branch_block_stmt_38/forx_xend273_bbx_xnph_PhiReq/$entry
      -- CP-element group 417: 	 branch_block_stmt_38/forx_xend273_bbx_xnph_PhiReq/$exit
      -- CP-element group 417: 	 branch_block_stmt_38/merge_stmt_1317_PhiReqMerge
      -- CP-element group 417: 	 branch_block_stmt_38/merge_stmt_1317_PhiAck/$entry
      -- CP-element group 417: 	 branch_block_stmt_38/merge_stmt_1317_PhiAck/$exit
      -- CP-element group 417: 	 branch_block_stmt_38/merge_stmt_1317_PhiAck/dummy
      -- 
    if_choice_transition_3076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1311_branch_ack_1, ack => convTranspose_CP_34_elements(417)); -- 
    cr_3098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(417), ack => type_cast_1338_inst_req_1); -- 
    rr_3093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(417), ack => type_cast_1338_inst_req_0); -- 
    -- CP-element group 418:  transition  place  input  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	416 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	496 
    -- CP-element group 418:  members (5) 
      -- CP-element group 418: 	 branch_block_stmt_38/forx_xend273_forx_xend500
      -- CP-element group 418: 	 branch_block_stmt_38/if_stmt_1311_else_link/else_choice_transition
      -- CP-element group 418: 	 branch_block_stmt_38/if_stmt_1311_else_link/$exit
      -- CP-element group 418: 	 branch_block_stmt_38/forx_xend273_forx_xend500_PhiReq/$entry
      -- CP-element group 418: 	 branch_block_stmt_38/forx_xend273_forx_xend500_PhiReq/$exit
      -- 
    else_choice_transition_3080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1311_branch_ack_0, ack => convTranspose_CP_34_elements(418)); -- 
    -- CP-element group 419:  transition  input  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	417 
    -- CP-element group 419: successors 
    -- CP-element group 419:  members (3) 
      -- CP-element group 419: 	 branch_block_stmt_38/assign_stmt_1323_to_assign_stmt_1352/type_cast_1338_Sample/ra
      -- CP-element group 419: 	 branch_block_stmt_38/assign_stmt_1323_to_assign_stmt_1352/type_cast_1338_Sample/$exit
      -- CP-element group 419: 	 branch_block_stmt_38/assign_stmt_1323_to_assign_stmt_1352/type_cast_1338_sample_completed_
      -- 
    ra_3094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1338_inst_ack_0, ack => convTranspose_CP_34_elements(419)); -- 
    -- CP-element group 420:  transition  place  input  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	417 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	490 
    -- CP-element group 420:  members (9) 
      -- CP-element group 420: 	 branch_block_stmt_38/assign_stmt_1323_to_assign_stmt_1352__exit__
      -- CP-element group 420: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427
      -- CP-element group 420: 	 branch_block_stmt_38/assign_stmt_1323_to_assign_stmt_1352/type_cast_1338_Update/ca
      -- CP-element group 420: 	 branch_block_stmt_38/assign_stmt_1323_to_assign_stmt_1352/type_cast_1338_Update/$exit
      -- CP-element group 420: 	 branch_block_stmt_38/assign_stmt_1323_to_assign_stmt_1352/type_cast_1338_update_completed_
      -- CP-element group 420: 	 branch_block_stmt_38/assign_stmt_1323_to_assign_stmt_1352/$exit
      -- CP-element group 420: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/$entry
      -- CP-element group 420: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1355/$entry
      -- CP-element group 420: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_sources/$entry
      -- 
    ca_3099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1338_inst_ack_1, ack => convTranspose_CP_34_elements(420)); -- 
    -- CP-element group 421:  transition  input  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	495 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	466 
    -- CP-element group 421:  members (3) 
      -- CP-element group 421: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_final_index_sum_regn_sample_complete
      -- CP-element group 421: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_final_index_sum_regn_Sample/$exit
      -- CP-element group 421: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_final_index_sum_regn_Sample/ack
      -- 
    ack_3128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1367_index_offset_ack_0, ack => convTranspose_CP_34_elements(421)); -- 
    -- CP-element group 422:  transition  input  output  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	495 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	423 
    -- CP-element group 422:  members (11) 
      -- CP-element group 422: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/addr_of_1368_sample_start_
      -- CP-element group 422: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_root_address_calculated
      -- CP-element group 422: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_offset_calculated
      -- CP-element group 422: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/addr_of_1368_request/req
      -- CP-element group 422: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/addr_of_1368_request/$entry
      -- CP-element group 422: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_base_plus_offset/sum_rename_ack
      -- CP-element group 422: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_base_plus_offset/sum_rename_req
      -- CP-element group 422: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_base_plus_offset/$exit
      -- CP-element group 422: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_base_plus_offset/$entry
      -- CP-element group 422: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_final_index_sum_regn_Update/ack
      -- CP-element group 422: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_final_index_sum_regn_Update/$exit
      -- 
    ack_3133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 422_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1367_index_offset_ack_1, ack => convTranspose_CP_34_elements(422)); -- 
    req_3142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(422), ack => addr_of_1368_final_reg_req_0); -- 
    -- CP-element group 423:  transition  input  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	422 
    -- CP-element group 423: successors 
    -- CP-element group 423:  members (3) 
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/addr_of_1368_sample_completed_
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/addr_of_1368_request/ack
      -- CP-element group 423: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/addr_of_1368_request/$exit
      -- 
    ack_3143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1368_final_reg_ack_0, ack => convTranspose_CP_34_elements(423)); -- 
    -- CP-element group 424:  join  fork  transition  input  output  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	495 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	425 
    -- CP-element group 424:  members (24) 
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/addr_of_1368_update_completed_
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Sample/word_access_start/word_0/rr
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Sample/word_access_start/word_0/$entry
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Sample/word_access_start/$entry
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_word_addrgen/root_register_ack
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_word_addrgen/root_register_req
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_word_addrgen/$exit
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_word_addrgen/$entry
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_base_plus_offset/sum_rename_ack
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_base_plus_offset/sum_rename_req
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_base_plus_offset/$exit
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_base_plus_offset/$entry
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_base_addr_resize/base_resize_ack
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_base_addr_resize/base_resize_req
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_base_addr_resize/$exit
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_base_addr_resize/$entry
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_base_address_resized
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_root_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_word_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_base_address_calculated
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_sample_start_
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/addr_of_1368_complete/ack
      -- CP-element group 424: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/addr_of_1368_complete/$exit
      -- 
    ack_3148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1368_final_reg_ack_1, ack => convTranspose_CP_34_elements(424)); -- 
    rr_3181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(424), ack => ptr_deref_1372_load_0_req_0); -- 
    -- CP-element group 425:  transition  input  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	424 
    -- CP-element group 425: successors 
    -- CP-element group 425:  members (5) 
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Sample/word_access_start/word_0/ra
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Sample/word_access_start/word_0/$exit
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Sample/word_access_start/$exit
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Sample/$exit
      -- CP-element group 425: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_sample_completed_
      -- 
    ra_3182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1372_load_0_ack_0, ack => convTranspose_CP_34_elements(425)); -- 
    -- CP-element group 426:  fork  transition  input  output  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	495 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	427 
    -- CP-element group 426: 	429 
    -- CP-element group 426: 	431 
    -- CP-element group 426: 	433 
    -- CP-element group 426: 	435 
    -- CP-element group 426: 	437 
    -- CP-element group 426: 	439 
    -- CP-element group 426: 	441 
    -- CP-element group 426:  members (33) 
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1426_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1426_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1396_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1376_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Update/ptr_deref_1372_Merge/merge_ack
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Update/word_access_complete/word_0/ca
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Update/ptr_deref_1372_Merge/merge_req
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1436_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1376_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Update/ptr_deref_1372_Merge/$entry
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1446_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1406_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Update/ptr_deref_1372_Merge/$exit
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1396_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1436_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1446_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Update/word_access_complete/word_0/$exit
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Update/word_access_complete/$exit
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1396_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1426_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Update/$exit
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1386_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1446_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1386_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1416_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1386_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1416_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1416_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_update_completed_
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1376_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1406_Sample/rr
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1406_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1436_Sample/rr
      -- 
    ca_3193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1372_load_0_ack_1, ack => convTranspose_CP_34_elements(426)); -- 
    rr_3206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(426), ack => type_cast_1376_inst_req_0); -- 
    rr_3220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(426), ack => type_cast_1386_inst_req_0); -- 
    rr_3234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(426), ack => type_cast_1396_inst_req_0); -- 
    rr_3248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(426), ack => type_cast_1406_inst_req_0); -- 
    rr_3262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(426), ack => type_cast_1416_inst_req_0); -- 
    rr_3276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(426), ack => type_cast_1426_inst_req_0); -- 
    rr_3290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(426), ack => type_cast_1436_inst_req_0); -- 
    rr_3304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(426), ack => type_cast_1446_inst_req_0); -- 
    -- CP-element group 427:  transition  input  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	426 
    -- CP-element group 427: successors 
    -- CP-element group 427:  members (3) 
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1376_sample_completed_
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1376_Sample/ra
      -- CP-element group 427: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1376_Sample/$exit
      -- 
    ra_3207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1376_inst_ack_0, ack => convTranspose_CP_34_elements(427)); -- 
    -- CP-element group 428:  transition  input  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	495 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	463 
    -- CP-element group 428:  members (3) 
      -- CP-element group 428: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1376_update_completed_
      -- CP-element group 428: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1376_Update/ca
      -- CP-element group 428: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1376_Update/$exit
      -- 
    ca_3212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1376_inst_ack_1, ack => convTranspose_CP_34_elements(428)); -- 
    -- CP-element group 429:  transition  input  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	426 
    -- CP-element group 429: successors 
    -- CP-element group 429:  members (3) 
      -- CP-element group 429: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1386_Sample/ra
      -- CP-element group 429: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1386_Sample/$exit
      -- CP-element group 429: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1386_sample_completed_
      -- 
    ra_3221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1386_inst_ack_0, ack => convTranspose_CP_34_elements(429)); -- 
    -- CP-element group 430:  transition  input  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	495 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	460 
    -- CP-element group 430:  members (3) 
      -- CP-element group 430: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1386_Update/ca
      -- CP-element group 430: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1386_Update/$exit
      -- CP-element group 430: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1386_update_completed_
      -- 
    ca_3226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1386_inst_ack_1, ack => convTranspose_CP_34_elements(430)); -- 
    -- CP-element group 431:  transition  input  bypass 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	426 
    -- CP-element group 431: successors 
    -- CP-element group 431:  members (3) 
      -- CP-element group 431: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1396_Sample/ra
      -- CP-element group 431: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1396_Sample/$exit
      -- CP-element group 431: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1396_sample_completed_
      -- 
    ra_3235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1396_inst_ack_0, ack => convTranspose_CP_34_elements(431)); -- 
    -- CP-element group 432:  transition  input  bypass 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	495 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	457 
    -- CP-element group 432:  members (3) 
      -- CP-element group 432: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1396_Update/$exit
      -- CP-element group 432: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1396_Update/ca
      -- CP-element group 432: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1396_update_completed_
      -- 
    ca_3240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1396_inst_ack_1, ack => convTranspose_CP_34_elements(432)); -- 
    -- CP-element group 433:  transition  input  bypass 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	426 
    -- CP-element group 433: successors 
    -- CP-element group 433:  members (3) 
      -- CP-element group 433: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1406_sample_completed_
      -- CP-element group 433: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1406_Sample/ra
      -- CP-element group 433: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1406_Sample/$exit
      -- 
    ra_3249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1406_inst_ack_0, ack => convTranspose_CP_34_elements(433)); -- 
    -- CP-element group 434:  transition  input  bypass 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	495 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	454 
    -- CP-element group 434:  members (3) 
      -- CP-element group 434: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1406_Update/ca
      -- CP-element group 434: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1406_Update/$exit
      -- CP-element group 434: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1406_update_completed_
      -- 
    ca_3254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 434_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1406_inst_ack_1, ack => convTranspose_CP_34_elements(434)); -- 
    -- CP-element group 435:  transition  input  bypass 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	426 
    -- CP-element group 435: successors 
    -- CP-element group 435:  members (3) 
      -- CP-element group 435: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1416_Sample/ra
      -- CP-element group 435: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1416_Sample/$exit
      -- CP-element group 435: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1416_sample_completed_
      -- 
    ra_3263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1416_inst_ack_0, ack => convTranspose_CP_34_elements(435)); -- 
    -- CP-element group 436:  transition  input  bypass 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	495 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	451 
    -- CP-element group 436:  members (3) 
      -- CP-element group 436: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1416_Update/ca
      -- CP-element group 436: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1416_Update/$exit
      -- CP-element group 436: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1416_update_completed_
      -- 
    ca_3268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1416_inst_ack_1, ack => convTranspose_CP_34_elements(436)); -- 
    -- CP-element group 437:  transition  input  bypass 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	426 
    -- CP-element group 437: successors 
    -- CP-element group 437:  members (3) 
      -- CP-element group 437: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1426_Sample/ra
      -- CP-element group 437: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1426_Sample/$exit
      -- CP-element group 437: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1426_sample_completed_
      -- 
    ra_3277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 437_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1426_inst_ack_0, ack => convTranspose_CP_34_elements(437)); -- 
    -- CP-element group 438:  transition  input  bypass 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	495 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	448 
    -- CP-element group 438:  members (3) 
      -- CP-element group 438: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1426_Update/$exit
      -- CP-element group 438: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1426_Update/ca
      -- CP-element group 438: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1426_update_completed_
      -- 
    ca_3282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 438_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1426_inst_ack_1, ack => convTranspose_CP_34_elements(438)); -- 
    -- CP-element group 439:  transition  input  bypass 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	426 
    -- CP-element group 439: successors 
    -- CP-element group 439:  members (3) 
      -- CP-element group 439: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1436_Sample/ra
      -- CP-element group 439: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1436_Sample/$exit
      -- CP-element group 439: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1436_sample_completed_
      -- 
    ra_3291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1436_inst_ack_0, ack => convTranspose_CP_34_elements(439)); -- 
    -- CP-element group 440:  transition  input  bypass 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	495 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	445 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1436_update_completed_
      -- CP-element group 440: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1436_Update/ca
      -- CP-element group 440: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1436_Update/$exit
      -- 
    ca_3296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1436_inst_ack_1, ack => convTranspose_CP_34_elements(440)); -- 
    -- CP-element group 441:  transition  input  bypass 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	426 
    -- CP-element group 441: successors 
    -- CP-element group 441:  members (3) 
      -- CP-element group 441: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1446_Sample/$exit
      -- CP-element group 441: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1446_sample_completed_
      -- CP-element group 441: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1446_Sample/ra
      -- 
    ra_3305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1446_inst_ack_0, ack => convTranspose_CP_34_elements(441)); -- 
    -- CP-element group 442:  transition  input  output  bypass 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	495 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	443 
    -- CP-element group 442:  members (6) 
      -- CP-element group 442: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1446_update_completed_
      -- CP-element group 442: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1448_Sample/req
      -- CP-element group 442: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1448_Sample/$entry
      -- CP-element group 442: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1448_sample_start_
      -- CP-element group 442: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1446_Update/ca
      -- CP-element group 442: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1446_Update/$exit
      -- 
    ca_3310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 442_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1446_inst_ack_1, ack => convTranspose_CP_34_elements(442)); -- 
    req_3318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(442), ack => WPIPE_ConvTranspose_output_pipe_1448_inst_req_0); -- 
    -- CP-element group 443:  transition  input  output  bypass 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	442 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	444 
    -- CP-element group 443:  members (6) 
      -- CP-element group 443: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1448_Update/req
      -- CP-element group 443: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1448_Update/$entry
      -- CP-element group 443: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1448_Sample/ack
      -- CP-element group 443: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1448_Sample/$exit
      -- CP-element group 443: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1448_update_start_
      -- CP-element group 443: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1448_sample_completed_
      -- 
    ack_3319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1448_inst_ack_0, ack => convTranspose_CP_34_elements(443)); -- 
    req_3323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(443), ack => WPIPE_ConvTranspose_output_pipe_1448_inst_req_1); -- 
    -- CP-element group 444:  transition  input  bypass 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	443 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	445 
    -- CP-element group 444:  members (3) 
      -- CP-element group 444: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1448_Update/ack
      -- CP-element group 444: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1448_Update/$exit
      -- CP-element group 444: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1448_update_completed_
      -- 
    ack_3324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1448_inst_ack_1, ack => convTranspose_CP_34_elements(444)); -- 
    -- CP-element group 445:  join  transition  output  bypass 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	440 
    -- CP-element group 445: 	444 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	446 
    -- CP-element group 445:  members (3) 
      -- CP-element group 445: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1451_Sample/req
      -- CP-element group 445: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1451_Sample/$entry
      -- CP-element group 445: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1451_sample_start_
      -- 
    req_3332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(445), ack => WPIPE_ConvTranspose_output_pipe_1451_inst_req_0); -- 
    convTranspose_cp_element_group_445: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_445"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(440) & convTranspose_CP_34_elements(444);
      gj_convTranspose_cp_element_group_445 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(445), clk => clk, reset => reset); --
    end block;
    -- CP-element group 446:  transition  input  output  bypass 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	445 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	447 
    -- CP-element group 446:  members (6) 
      -- CP-element group 446: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1451_Update/req
      -- CP-element group 446: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1451_Update/$entry
      -- CP-element group 446: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1451_Sample/ack
      -- CP-element group 446: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1451_Sample/$exit
      -- CP-element group 446: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1451_update_start_
      -- CP-element group 446: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1451_sample_completed_
      -- 
    ack_3333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 446_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1451_inst_ack_0, ack => convTranspose_CP_34_elements(446)); -- 
    req_3337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(446), ack => WPIPE_ConvTranspose_output_pipe_1451_inst_req_1); -- 
    -- CP-element group 447:  transition  input  bypass 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	446 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	448 
    -- CP-element group 447:  members (3) 
      -- CP-element group 447: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1451_Update/ack
      -- CP-element group 447: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1451_Update/$exit
      -- CP-element group 447: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1451_update_completed_
      -- 
    ack_3338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1451_inst_ack_1, ack => convTranspose_CP_34_elements(447)); -- 
    -- CP-element group 448:  join  transition  output  bypass 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	438 
    -- CP-element group 448: 	447 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	449 
    -- CP-element group 448:  members (3) 
      -- CP-element group 448: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1454_sample_start_
      -- CP-element group 448: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1454_Sample/req
      -- CP-element group 448: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1454_Sample/$entry
      -- 
    req_3346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(448), ack => WPIPE_ConvTranspose_output_pipe_1454_inst_req_0); -- 
    convTranspose_cp_element_group_448: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_448"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(438) & convTranspose_CP_34_elements(447);
      gj_convTranspose_cp_element_group_448 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(448), clk => clk, reset => reset); --
    end block;
    -- CP-element group 449:  transition  input  output  bypass 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	448 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	450 
    -- CP-element group 449:  members (6) 
      -- CP-element group 449: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1454_sample_completed_
      -- CP-element group 449: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1454_Update/req
      -- CP-element group 449: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1454_Update/$entry
      -- CP-element group 449: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1454_Sample/ack
      -- CP-element group 449: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1454_Sample/$exit
      -- CP-element group 449: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1454_update_start_
      -- 
    ack_3347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 449_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1454_inst_ack_0, ack => convTranspose_CP_34_elements(449)); -- 
    req_3351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(449), ack => WPIPE_ConvTranspose_output_pipe_1454_inst_req_1); -- 
    -- CP-element group 450:  transition  input  bypass 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	449 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	451 
    -- CP-element group 450:  members (3) 
      -- CP-element group 450: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1454_Update/ack
      -- CP-element group 450: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1454_Update/$exit
      -- CP-element group 450: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1454_update_completed_
      -- 
    ack_3352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 450_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1454_inst_ack_1, ack => convTranspose_CP_34_elements(450)); -- 
    -- CP-element group 451:  join  transition  output  bypass 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	436 
    -- CP-element group 451: 	450 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	452 
    -- CP-element group 451:  members (3) 
      -- CP-element group 451: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1457_Sample/req
      -- CP-element group 451: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1457_Sample/$entry
      -- CP-element group 451: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1457_sample_start_
      -- 
    req_3360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(451), ack => WPIPE_ConvTranspose_output_pipe_1457_inst_req_0); -- 
    convTranspose_cp_element_group_451: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_451"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(436) & convTranspose_CP_34_elements(450);
      gj_convTranspose_cp_element_group_451 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(451), clk => clk, reset => reset); --
    end block;
    -- CP-element group 452:  transition  input  output  bypass 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	451 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	453 
    -- CP-element group 452:  members (6) 
      -- CP-element group 452: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1457_Update/req
      -- CP-element group 452: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1457_Update/$entry
      -- CP-element group 452: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1457_Sample/ack
      -- CP-element group 452: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1457_Sample/$exit
      -- CP-element group 452: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1457_update_start_
      -- CP-element group 452: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1457_sample_completed_
      -- 
    ack_3361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 452_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1457_inst_ack_0, ack => convTranspose_CP_34_elements(452)); -- 
    req_3365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(452), ack => WPIPE_ConvTranspose_output_pipe_1457_inst_req_1); -- 
    -- CP-element group 453:  transition  input  bypass 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	452 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	454 
    -- CP-element group 453:  members (3) 
      -- CP-element group 453: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1457_Update/ack
      -- CP-element group 453: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1457_Update/$exit
      -- CP-element group 453: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1457_update_completed_
      -- 
    ack_3366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1457_inst_ack_1, ack => convTranspose_CP_34_elements(453)); -- 
    -- CP-element group 454:  join  transition  output  bypass 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	434 
    -- CP-element group 454: 	453 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	455 
    -- CP-element group 454:  members (3) 
      -- CP-element group 454: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1460_Sample/req
      -- CP-element group 454: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1460_Sample/$entry
      -- CP-element group 454: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1460_sample_start_
      -- 
    req_3374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(454), ack => WPIPE_ConvTranspose_output_pipe_1460_inst_req_0); -- 
    convTranspose_cp_element_group_454: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_454"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(434) & convTranspose_CP_34_elements(453);
      gj_convTranspose_cp_element_group_454 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(454), clk => clk, reset => reset); --
    end block;
    -- CP-element group 455:  transition  input  output  bypass 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	454 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	456 
    -- CP-element group 455:  members (6) 
      -- CP-element group 455: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1460_Sample/ack
      -- CP-element group 455: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1460_Sample/$exit
      -- CP-element group 455: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1460_update_start_
      -- CP-element group 455: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1460_sample_completed_
      -- CP-element group 455: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1460_Update/$entry
      -- CP-element group 455: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1460_Update/req
      -- 
    ack_3375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 455_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1460_inst_ack_0, ack => convTranspose_CP_34_elements(455)); -- 
    req_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(455), ack => WPIPE_ConvTranspose_output_pipe_1460_inst_req_1); -- 
    -- CP-element group 456:  transition  input  bypass 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	455 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	457 
    -- CP-element group 456:  members (3) 
      -- CP-element group 456: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1460_update_completed_
      -- CP-element group 456: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1460_Update/$exit
      -- CP-element group 456: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1460_Update/ack
      -- 
    ack_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 456_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1460_inst_ack_1, ack => convTranspose_CP_34_elements(456)); -- 
    -- CP-element group 457:  join  transition  output  bypass 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	432 
    -- CP-element group 457: 	456 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	458 
    -- CP-element group 457:  members (3) 
      -- CP-element group 457: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1463_sample_start_
      -- CP-element group 457: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1463_Sample/$entry
      -- CP-element group 457: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1463_Sample/req
      -- 
    req_3388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(457), ack => WPIPE_ConvTranspose_output_pipe_1463_inst_req_0); -- 
    convTranspose_cp_element_group_457: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_457"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(432) & convTranspose_CP_34_elements(456);
      gj_convTranspose_cp_element_group_457 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(457), clk => clk, reset => reset); --
    end block;
    -- CP-element group 458:  transition  input  output  bypass 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	457 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	459 
    -- CP-element group 458:  members (6) 
      -- CP-element group 458: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1463_sample_completed_
      -- CP-element group 458: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1463_update_start_
      -- CP-element group 458: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1463_Sample/$exit
      -- CP-element group 458: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1463_Sample/ack
      -- CP-element group 458: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1463_Update/$entry
      -- CP-element group 458: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1463_Update/req
      -- 
    ack_3389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 458_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1463_inst_ack_0, ack => convTranspose_CP_34_elements(458)); -- 
    req_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(458), ack => WPIPE_ConvTranspose_output_pipe_1463_inst_req_1); -- 
    -- CP-element group 459:  transition  input  bypass 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	458 
    -- CP-element group 459: successors 
    -- CP-element group 459: 	460 
    -- CP-element group 459:  members (3) 
      -- CP-element group 459: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1463_update_completed_
      -- CP-element group 459: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1463_Update/$exit
      -- CP-element group 459: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1463_Update/ack
      -- 
    ack_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 459_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1463_inst_ack_1, ack => convTranspose_CP_34_elements(459)); -- 
    -- CP-element group 460:  join  transition  output  bypass 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	430 
    -- CP-element group 460: 	459 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	461 
    -- CP-element group 460:  members (3) 
      -- CP-element group 460: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1466_sample_start_
      -- CP-element group 460: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1466_Sample/$entry
      -- CP-element group 460: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1466_Sample/req
      -- 
    req_3402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(460), ack => WPIPE_ConvTranspose_output_pipe_1466_inst_req_0); -- 
    convTranspose_cp_element_group_460: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_460"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(430) & convTranspose_CP_34_elements(459);
      gj_convTranspose_cp_element_group_460 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(460), clk => clk, reset => reset); --
    end block;
    -- CP-element group 461:  transition  input  output  bypass 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	460 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	462 
    -- CP-element group 461:  members (6) 
      -- CP-element group 461: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1466_sample_completed_
      -- CP-element group 461: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1466_update_start_
      -- CP-element group 461: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1466_Sample/$exit
      -- CP-element group 461: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1466_Sample/ack
      -- CP-element group 461: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1466_Update/$entry
      -- CP-element group 461: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1466_Update/req
      -- 
    ack_3403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 461_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1466_inst_ack_0, ack => convTranspose_CP_34_elements(461)); -- 
    req_3407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(461), ack => WPIPE_ConvTranspose_output_pipe_1466_inst_req_1); -- 
    -- CP-element group 462:  transition  input  bypass 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	461 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	463 
    -- CP-element group 462:  members (3) 
      -- CP-element group 462: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1466_update_completed_
      -- CP-element group 462: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1466_Update/$exit
      -- CP-element group 462: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1466_Update/ack
      -- 
    ack_3408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 462_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1466_inst_ack_1, ack => convTranspose_CP_34_elements(462)); -- 
    -- CP-element group 463:  join  transition  output  bypass 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	428 
    -- CP-element group 463: 	462 
    -- CP-element group 463: successors 
    -- CP-element group 463: 	464 
    -- CP-element group 463:  members (3) 
      -- CP-element group 463: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1469_sample_start_
      -- CP-element group 463: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1469_Sample/$entry
      -- CP-element group 463: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1469_Sample/req
      -- 
    req_3416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(463), ack => WPIPE_ConvTranspose_output_pipe_1469_inst_req_0); -- 
    convTranspose_cp_element_group_463: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_463"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(428) & convTranspose_CP_34_elements(462);
      gj_convTranspose_cp_element_group_463 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(463), clk => clk, reset => reset); --
    end block;
    -- CP-element group 464:  transition  input  output  bypass 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	463 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	465 
    -- CP-element group 464:  members (6) 
      -- CP-element group 464: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1469_sample_completed_
      -- CP-element group 464: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1469_update_start_
      -- CP-element group 464: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1469_Sample/$exit
      -- CP-element group 464: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1469_Sample/ack
      -- CP-element group 464: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1469_Update/$entry
      -- CP-element group 464: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1469_Update/req
      -- 
    ack_3417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 464_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1469_inst_ack_0, ack => convTranspose_CP_34_elements(464)); -- 
    req_3421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(464), ack => WPIPE_ConvTranspose_output_pipe_1469_inst_req_1); -- 
    -- CP-element group 465:  transition  input  bypass 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	464 
    -- CP-element group 465: successors 
    -- CP-element group 465: 	466 
    -- CP-element group 465:  members (3) 
      -- CP-element group 465: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1469_update_completed_
      -- CP-element group 465: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1469_Update/$exit
      -- CP-element group 465: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/WPIPE_ConvTranspose_output_pipe_1469_Update/ack
      -- 
    ack_3422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1469_inst_ack_1, ack => convTranspose_CP_34_elements(465)); -- 
    -- CP-element group 466:  branch  join  transition  place  output  bypass 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	421 
    -- CP-element group 466: 	465 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	467 
    -- CP-element group 466: 	468 
    -- CP-element group 466:  members (10) 
      -- CP-element group 466: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482__exit__
      -- CP-element group 466: 	 branch_block_stmt_38/if_stmt_1483__entry__
      -- CP-element group 466: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/$exit
      -- CP-element group 466: 	 branch_block_stmt_38/if_stmt_1483_dead_link/$entry
      -- CP-element group 466: 	 branch_block_stmt_38/if_stmt_1483_eval_test/$entry
      -- CP-element group 466: 	 branch_block_stmt_38/if_stmt_1483_eval_test/$exit
      -- CP-element group 466: 	 branch_block_stmt_38/if_stmt_1483_eval_test/branch_req
      -- CP-element group 466: 	 branch_block_stmt_38/R_exitcond1_1484_place
      -- CP-element group 466: 	 branch_block_stmt_38/if_stmt_1483_if_link/$entry
      -- CP-element group 466: 	 branch_block_stmt_38/if_stmt_1483_else_link/$entry
      -- 
    branch_req_3430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(466), ack => if_stmt_1483_branch_req_0); -- 
    convTranspose_cp_element_group_466: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_466"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(421) & convTranspose_CP_34_elements(465);
      gj_convTranspose_cp_element_group_466 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(466), clk => clk, reset => reset); --
    end block;
    -- CP-element group 467:  merge  transition  place  input  bypass 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	466 
    -- CP-element group 467: successors 
    -- CP-element group 467: 	496 
    -- CP-element group 467:  members (13) 
      -- CP-element group 467: 	 branch_block_stmt_38/merge_stmt_1489__exit__
      -- CP-element group 467: 	 branch_block_stmt_38/forx_xend500x_xloopexit_forx_xend500
      -- CP-element group 467: 	 branch_block_stmt_38/if_stmt_1483_if_link/$exit
      -- CP-element group 467: 	 branch_block_stmt_38/if_stmt_1483_if_link/if_choice_transition
      -- CP-element group 467: 	 branch_block_stmt_38/forx_xbody427_forx_xend500x_xloopexit
      -- CP-element group 467: 	 branch_block_stmt_38/forx_xbody427_forx_xend500x_xloopexit_PhiReq/$entry
      -- CP-element group 467: 	 branch_block_stmt_38/forx_xbody427_forx_xend500x_xloopexit_PhiReq/$exit
      -- CP-element group 467: 	 branch_block_stmt_38/merge_stmt_1489_PhiReqMerge
      -- CP-element group 467: 	 branch_block_stmt_38/merge_stmt_1489_PhiAck/$entry
      -- CP-element group 467: 	 branch_block_stmt_38/merge_stmt_1489_PhiAck/$exit
      -- CP-element group 467: 	 branch_block_stmt_38/merge_stmt_1489_PhiAck/dummy
      -- CP-element group 467: 	 branch_block_stmt_38/forx_xend500x_xloopexit_forx_xend500_PhiReq/$entry
      -- CP-element group 467: 	 branch_block_stmt_38/forx_xend500x_xloopexit_forx_xend500_PhiReq/$exit
      -- 
    if_choice_transition_3435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 467_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1483_branch_ack_1, ack => convTranspose_CP_34_elements(467)); -- 
    -- CP-element group 468:  fork  transition  place  input  output  bypass 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	466 
    -- CP-element group 468: successors 
    -- CP-element group 468: 	491 
    -- CP-element group 468: 	492 
    -- CP-element group 468:  members (12) 
      -- CP-element group 468: 	 branch_block_stmt_38/if_stmt_1483_else_link/$exit
      -- CP-element group 468: 	 branch_block_stmt_38/if_stmt_1483_else_link/else_choice_transition
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/$entry
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1355/$entry
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_sources/$entry
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_sources/type_cast_1361/$entry
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_sources/type_cast_1361/SplitProtocol/$entry
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_sources/type_cast_1361/SplitProtocol/Sample/$entry
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_sources/type_cast_1361/SplitProtocol/Sample/rr
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_sources/type_cast_1361/SplitProtocol/Update/$entry
      -- CP-element group 468: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_sources/type_cast_1361/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1483_branch_ack_0, ack => convTranspose_CP_34_elements(468)); -- 
    rr_3714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(468), ack => type_cast_1361_inst_req_0); -- 
    cr_3719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(468), ack => type_cast_1361_inst_req_1); -- 
    -- CP-element group 469:  merge  branch  transition  place  output  bypass 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	165 
    -- CP-element group 469: 	120 
    -- CP-element group 469: successors 
    -- CP-element group 469: 	121 
    -- CP-element group 469: 	122 
    -- CP-element group 469:  members (17) 
      -- CP-element group 469: 	 branch_block_stmt_38/merge_stmt_429__exit__
      -- CP-element group 469: 	 branch_block_stmt_38/assign_stmt_435__entry__
      -- CP-element group 469: 	 branch_block_stmt_38/assign_stmt_435__exit__
      -- CP-element group 469: 	 branch_block_stmt_38/if_stmt_436__entry__
      -- CP-element group 469: 	 branch_block_stmt_38/assign_stmt_435/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/assign_stmt_435/$exit
      -- CP-element group 469: 	 branch_block_stmt_38/if_stmt_436_dead_link/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/if_stmt_436_eval_test/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/if_stmt_436_eval_test/$exit
      -- CP-element group 469: 	 branch_block_stmt_38/if_stmt_436_eval_test/branch_req
      -- CP-element group 469: 	 branch_block_stmt_38/R_cmp194509_437_place
      -- CP-element group 469: 	 branch_block_stmt_38/if_stmt_436_if_link/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/if_stmt_436_else_link/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/merge_stmt_429_PhiReqMerge
      -- CP-element group 469: 	 branch_block_stmt_38/merge_stmt_429_PhiAck/$entry
      -- CP-element group 469: 	 branch_block_stmt_38/merge_stmt_429_PhiAck/$exit
      -- CP-element group 469: 	 branch_block_stmt_38/merge_stmt_429_PhiAck/dummy
      -- 
    branch_req_922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(469), ack => if_stmt_436_branch_req_0); -- 
    convTranspose_CP_34_elements(469) <= OrReduce(convTranspose_CP_34_elements(165) & convTranspose_CP_34_elements(120));
    -- CP-element group 470:  transition  output  delay-element  bypass 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	124 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	474 
    -- CP-element group 470:  members (5) 
      -- CP-element group 470: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/$exit
      -- CP-element group 470: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_474/$exit
      -- CP-element group 470: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/$exit
      -- CP-element group 470: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_478_konst_delay_trans
      -- CP-element group 470: 	 branch_block_stmt_38/bbx_xnph515_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_req
      -- 
    phi_stmt_474_req_3487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_474_req_3487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(470), ack => phi_stmt_474_req_0); -- 
    -- Element group convTranspose_CP_34_elements(470) is a control-delay.
    cp_element_470_delay: control_delay_element  generic map(name => " 470_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(124), ack => convTranspose_CP_34_elements(470), clk => clk, reset =>reset);
    -- CP-element group 471:  transition  input  bypass 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	166 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	473 
    -- CP-element group 471:  members (2) 
      -- CP-element group 471: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Sample/$exit
      -- CP-element group 471: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Sample/ra
      -- 
    ra_3507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 471_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_480_inst_ack_0, ack => convTranspose_CP_34_elements(471)); -- 
    -- CP-element group 472:  transition  input  bypass 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	166 
    -- CP-element group 472: successors 
    -- CP-element group 472: 	473 
    -- CP-element group 472:  members (2) 
      -- CP-element group 472: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Update/$exit
      -- CP-element group 472: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/Update/ca
      -- 
    ca_3512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 472_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_480_inst_ack_1, ack => convTranspose_CP_34_elements(472)); -- 
    -- CP-element group 473:  join  transition  output  bypass 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	471 
    -- CP-element group 473: 	472 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	474 
    -- CP-element group 473:  members (6) 
      -- CP-element group 473: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 473: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/$exit
      -- CP-element group 473: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/$exit
      -- CP-element group 473: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/$exit
      -- CP-element group 473: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_sources/type_cast_480/SplitProtocol/$exit
      -- CP-element group 473: 	 branch_block_stmt_38/forx_xbody_forx_xbody_PhiReq/phi_stmt_474/phi_stmt_474_req
      -- 
    phi_stmt_474_req_3513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_474_req_3513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(473), ack => phi_stmt_474_req_1); -- 
    convTranspose_cp_element_group_473: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_473"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(471) & convTranspose_CP_34_elements(472);
      gj_convTranspose_cp_element_group_473 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(473), clk => clk, reset => reset); --
    end block;
    -- CP-element group 474:  merge  transition  place  bypass 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	470 
    -- CP-element group 474: 	473 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	475 
    -- CP-element group 474:  members (2) 
      -- CP-element group 474: 	 branch_block_stmt_38/merge_stmt_473_PhiReqMerge
      -- CP-element group 474: 	 branch_block_stmt_38/merge_stmt_473_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(474) <= OrReduce(convTranspose_CP_34_elements(470) & convTranspose_CP_34_elements(473));
    -- CP-element group 475:  fork  transition  place  input  output  bypass 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	474 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	163 
    -- CP-element group 475: 	125 
    -- CP-element group 475: 	126 
    -- CP-element group 475: 	128 
    -- CP-element group 475: 	129 
    -- CP-element group 475: 	132 
    -- CP-element group 475: 	136 
    -- CP-element group 475: 	140 
    -- CP-element group 475: 	144 
    -- CP-element group 475: 	148 
    -- CP-element group 475: 	152 
    -- CP-element group 475: 	156 
    -- CP-element group 475: 	160 
    -- CP-element group 475:  members (56) 
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_update_start_
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_update_start_
      -- CP-element group 475: 	 branch_block_stmt_38/merge_stmt_473__exit__
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636__entry__
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_597_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_543_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/word_access_complete/word_0/cr
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/word_access_complete/word_0/$entry
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/word_access_complete/$entry
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_579_update_start_
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_615_update_start_
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_561_update_start_
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/ptr_deref_623_update_start_
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/$entry
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_update_start_
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_resized_1
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_scaled_1
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_computed_1
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_resize_1/$entry
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_resize_1/$exit
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_resize_1/index_resize_req
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_resize_1/index_resize_ack
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_scale_1/$entry
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_scale_1/$exit
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_scale_1/scale_rename_req
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_index_scale_1/scale_rename_ack
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_update_start
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Sample/$entry
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Sample/req
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/array_obj_ref_486_final_index_sum_regn_Update/req
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_complete/$entry
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/addr_of_487_complete/req
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_sample_start_
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Sample/$entry
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/RPIPE_ConvTranspose_input_pipe_490_Sample/rr
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_update_start_
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_494_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_update_start_
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_507_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_update_start_
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_38/assign_stmt_488_to_assign_stmt_636/type_cast_525_Update/cr
      -- CP-element group 475: 	 branch_block_stmt_38/merge_stmt_473_PhiAck/$exit
      -- CP-element group 475: 	 branch_block_stmt_38/merge_stmt_473_PhiAck/phi_stmt_474_ack
      -- 
    phi_stmt_474_ack_3518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 475_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_474_ack_0, ack => convTranspose_CP_34_elements(475)); -- 
    cr_1194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(475), ack => type_cast_597_inst_req_1); -- 
    cr_1110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(475), ack => type_cast_543_inst_req_1); -- 
    cr_1272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(475), ack => ptr_deref_623_store_0_req_1); -- 
    cr_1222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(475), ack => type_cast_615_inst_req_1); -- 
    cr_1166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(475), ack => type_cast_579_inst_req_1); -- 
    cr_1138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(475), ack => type_cast_561_inst_req_1); -- 
    req_978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(475), ack => array_obj_ref_486_index_offset_req_0); -- 
    req_983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(475), ack => array_obj_ref_486_index_offset_req_1); -- 
    req_998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(475), ack => addr_of_487_final_reg_req_1); -- 
    rr_1007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(475), ack => RPIPE_ConvTranspose_input_pipe_490_inst_req_0); -- 
    cr_1026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(475), ack => type_cast_494_inst_req_1); -- 
    cr_1054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(475), ack => type_cast_507_inst_req_1); -- 
    cr_1082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(475), ack => type_cast_525_inst_req_1); -- 
    -- CP-element group 476:  transition  output  delay-element  bypass 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	168 
    -- CP-element group 476: successors 
    -- CP-element group 476: 	480 
    -- CP-element group 476:  members (5) 
      -- CP-element group 476: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/$exit
      -- CP-element group 476: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_681/$exit
      -- CP-element group 476: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/$exit
      -- CP-element group 476: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_685_konst_delay_trans
      -- CP-element group 476: 	 branch_block_stmt_38/bbx_xnph511_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_req
      -- 
    phi_stmt_681_req_3541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_681_req_3541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(476), ack => phi_stmt_681_req_0); -- 
    -- Element group convTranspose_CP_34_elements(476) is a control-delay.
    cp_element_476_delay: control_delay_element  generic map(name => " 476_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(168), ack => convTranspose_CP_34_elements(476), clk => clk, reset =>reset);
    -- CP-element group 477:  transition  input  bypass 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	210 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	479 
    -- CP-element group 477:  members (2) 
      -- CP-element group 477: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Sample/$exit
      -- CP-element group 477: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Sample/ra
      -- 
    ra_3561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 477_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_687_inst_ack_0, ack => convTranspose_CP_34_elements(477)); -- 
    -- CP-element group 478:  transition  input  bypass 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	210 
    -- CP-element group 478: successors 
    -- CP-element group 478: 	479 
    -- CP-element group 478:  members (2) 
      -- CP-element group 478: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Update/$exit
      -- CP-element group 478: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/Update/ca
      -- 
    ca_3566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 478_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_687_inst_ack_1, ack => convTranspose_CP_34_elements(478)); -- 
    -- CP-element group 479:  join  transition  output  bypass 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	477 
    -- CP-element group 479: 	478 
    -- CP-element group 479: successors 
    -- CP-element group 479: 	480 
    -- CP-element group 479:  members (6) 
      -- CP-element group 479: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/$exit
      -- CP-element group 479: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/$exit
      -- CP-element group 479: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/$exit
      -- CP-element group 479: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/$exit
      -- CP-element group 479: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_sources/type_cast_687/SplitProtocol/$exit
      -- CP-element group 479: 	 branch_block_stmt_38/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_681/phi_stmt_681_req
      -- 
    phi_stmt_681_req_3567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_681_req_3567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(479), ack => phi_stmt_681_req_1); -- 
    convTranspose_cp_element_group_479: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_479"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(477) & convTranspose_CP_34_elements(478);
      gj_convTranspose_cp_element_group_479 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(479), clk => clk, reset => reset); --
    end block;
    -- CP-element group 480:  merge  transition  place  bypass 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	476 
    -- CP-element group 480: 	479 
    -- CP-element group 480: successors 
    -- CP-element group 480: 	481 
    -- CP-element group 480:  members (2) 
      -- CP-element group 480: 	 branch_block_stmt_38/merge_stmt_680_PhiReqMerge
      -- CP-element group 480: 	 branch_block_stmt_38/merge_stmt_680_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(480) <= OrReduce(convTranspose_CP_34_elements(476) & convTranspose_CP_34_elements(479));
    -- CP-element group 481:  fork  transition  place  input  output  bypass 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	480 
    -- CP-element group 481: successors 
    -- CP-element group 481: 	180 
    -- CP-element group 481: 	184 
    -- CP-element group 481: 	188 
    -- CP-element group 481: 	172 
    -- CP-element group 481: 	173 
    -- CP-element group 481: 	176 
    -- CP-element group 481: 	192 
    -- CP-element group 481: 	196 
    -- CP-element group 481: 	200 
    -- CP-element group 481: 	204 
    -- CP-element group 481: 	207 
    -- CP-element group 481: 	169 
    -- CP-element group 481: 	170 
    -- CP-element group 481:  members (56) 
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_update_start_
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_update_start_
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_update_start_
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Sample/$entry
      -- CP-element group 481: 	 branch_block_stmt_38/merge_stmt_680__exit__
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843__entry__
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_update_start_
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_complete/req
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/$entry
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_complete/$entry
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/addr_of_694_update_start_
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Update/req
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_sample_start_
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Sample/req
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/RPIPE_ConvTranspose_input_pipe_697_Sample/rr
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_Sample/$entry
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_714_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_732_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_resized_1
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_final_index_sum_regn_update_start
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_scale_1/scale_rename_ack
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_scale_1/scale_rename_req
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_scale_1/$exit
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_scale_1/$entry
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_resize_1/index_resize_ack
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_resize_1/index_resize_req
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_701_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_resize_1/$exit
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_resize_1/$entry
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_computed_1
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/array_obj_ref_693_index_scaled_1
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_750_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_update_start_
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_768_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_update_start_
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_786_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_update_start_
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_804_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_update_start_
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/type_cast_822_Update/cr
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_update_start_
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/$entry
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/word_access_complete/$entry
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/word_access_complete/word_0/$entry
      -- CP-element group 481: 	 branch_block_stmt_38/assign_stmt_695_to_assign_stmt_843/ptr_deref_830_Update/word_access_complete/word_0/cr
      -- CP-element group 481: 	 branch_block_stmt_38/merge_stmt_680_PhiAck/$exit
      -- CP-element group 481: 	 branch_block_stmt_38/merge_stmt_680_PhiAck/phi_stmt_681_ack
      -- 
    phi_stmt_681_ack_3572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 481_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_681_ack_0, ack => convTranspose_CP_34_elements(481)); -- 
    req_1357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(481), ack => addr_of_694_final_reg_req_1); -- 
    req_1342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(481), ack => array_obj_ref_693_index_offset_req_1); -- 
    req_1337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(481), ack => array_obj_ref_693_index_offset_req_0); -- 
    cr_1441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(481), ack => type_cast_732_inst_req_1); -- 
    rr_1366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(481), ack => RPIPE_ConvTranspose_input_pipe_697_inst_req_0); -- 
    cr_1413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(481), ack => type_cast_714_inst_req_1); -- 
    cr_1385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(481), ack => type_cast_701_inst_req_1); -- 
    cr_1469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(481), ack => type_cast_750_inst_req_1); -- 
    cr_1497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(481), ack => type_cast_768_inst_req_1); -- 
    cr_1525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(481), ack => type_cast_786_inst_req_1); -- 
    cr_1553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(481), ack => type_cast_804_inst_req_1); -- 
    cr_1581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(481), ack => type_cast_822_inst_req_1); -- 
    cr_1631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(481), ack => ptr_deref_830_store_0_req_1); -- 
    -- CP-element group 482:  merge  fork  transition  place  output  bypass 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	209 
    -- CP-element group 482: 	122 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	211 
    -- CP-element group 482: 	212 
    -- CP-element group 482: 	213 
    -- CP-element group 482: 	214 
    -- CP-element group 482: 	215 
    -- CP-element group 482: 	216 
    -- CP-element group 482:  members (25) 
      -- CP-element group 482: 	 branch_block_stmt_38/merge_stmt_852__exit__
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880__entry__
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Sample/rr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_855_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Sample/rr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_859_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_update_start_
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Sample/rr
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/assign_stmt_856_to_assign_stmt_880/type_cast_863_Update/cr
      -- CP-element group 482: 	 branch_block_stmt_38/merge_stmt_852_PhiReqMerge
      -- CP-element group 482: 	 branch_block_stmt_38/merge_stmt_852_PhiAck/$entry
      -- CP-element group 482: 	 branch_block_stmt_38/merge_stmt_852_PhiAck/$exit
      -- CP-element group 482: 	 branch_block_stmt_38/merge_stmt_852_PhiAck/dummy
      -- 
    rr_1662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_855_inst_req_0); -- 
    cr_1667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_855_inst_req_1); -- 
    rr_1676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_859_inst_req_0); -- 
    cr_1681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_859_inst_req_1); -- 
    rr_1690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_863_inst_req_0); -- 
    cr_1695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(482), ack => type_cast_863_inst_req_1); -- 
    convTranspose_CP_34_elements(482) <= OrReduce(convTranspose_CP_34_elements(209) & convTranspose_CP_34_elements(122));
    -- CP-element group 483:  transition  output  delay-element  bypass 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	221 
    -- CP-element group 483: successors 
    -- CP-element group 483: 	487 
    -- CP-element group 483:  members (5) 
      -- CP-element group 483: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/$exit
      -- CP-element group 483: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_925/$exit
      -- CP-element group 483: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/$exit
      -- CP-element group 483: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_931_konst_delay_trans
      -- CP-element group 483: 	 branch_block_stmt_38/bbx_xnph507_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_req
      -- 
    phi_stmt_925_req_3618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_925_req_3618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(483), ack => phi_stmt_925_req_1); -- 
    -- Element group convTranspose_CP_34_elements(483) is a control-delay.
    cp_element_483_delay: control_delay_element  generic map(name => " 483_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(221), ack => convTranspose_CP_34_elements(483), clk => clk, reset =>reset);
    -- CP-element group 484:  transition  input  bypass 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	230 
    -- CP-element group 484: successors 
    -- CP-element group 484: 	486 
    -- CP-element group 484:  members (2) 
      -- CP-element group 484: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Sample/$exit
      -- CP-element group 484: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Sample/ra
      -- 
    ra_3638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 484_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_928_inst_ack_0, ack => convTranspose_CP_34_elements(484)); -- 
    -- CP-element group 485:  transition  input  bypass 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	230 
    -- CP-element group 485: successors 
    -- CP-element group 485: 	486 
    -- CP-element group 485:  members (2) 
      -- CP-element group 485: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Update/$exit
      -- CP-element group 485: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/Update/ca
      -- 
    ca_3643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_928_inst_ack_1, ack => convTranspose_CP_34_elements(485)); -- 
    -- CP-element group 486:  join  transition  output  bypass 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	484 
    -- CP-element group 486: 	485 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	487 
    -- CP-element group 486:  members (6) 
      -- CP-element group 486: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/$exit
      -- CP-element group 486: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/$exit
      -- CP-element group 486: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/$exit
      -- CP-element group 486: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/$exit
      -- CP-element group 486: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_sources/type_cast_928/SplitProtocol/$exit
      -- CP-element group 486: 	 branch_block_stmt_38/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_925/phi_stmt_925_req
      -- 
    phi_stmt_925_req_3644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_925_req_3644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(486), ack => phi_stmt_925_req_0); -- 
    convTranspose_cp_element_group_486: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_486"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(484) & convTranspose_CP_34_elements(485);
      gj_convTranspose_cp_element_group_486 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(486), clk => clk, reset => reset); --
    end block;
    -- CP-element group 487:  merge  transition  place  bypass 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	483 
    -- CP-element group 487: 	486 
    -- CP-element group 487: successors 
    -- CP-element group 487: 	488 
    -- CP-element group 487:  members (2) 
      -- CP-element group 487: 	 branch_block_stmt_38/merge_stmt_924_PhiReqMerge
      -- CP-element group 487: 	 branch_block_stmt_38/merge_stmt_924_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(487) <= OrReduce(convTranspose_CP_34_elements(483) & convTranspose_CP_34_elements(486));
    -- CP-element group 488:  fork  transition  place  input  output  bypass 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	487 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	222 
    -- CP-element group 488: 	223 
    -- CP-element group 488: 	225 
    -- CP-element group 488: 	227 
    -- CP-element group 488:  members (29) 
      -- CP-element group 488: 	 branch_block_stmt_38/merge_stmt_924__exit__
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955__entry__
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/$entry
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_update_start_
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_resized_1
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_scaled_1
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_computed_1
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_resize_1/$entry
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_resize_1/$exit
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_resize_1/index_resize_req
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_resize_1/index_resize_ack
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_scale_1/$entry
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_scale_1/$exit
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_scale_1/scale_rename_req
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_index_scale_1/scale_rename_ack
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_update_start
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Sample/$entry
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Sample/req
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Update/$entry
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/array_obj_ref_937_final_index_sum_regn_Update/req
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_complete/$entry
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/addr_of_938_complete/req
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_update_start_
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/$entry
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/word_access_complete/$entry
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/word_access_complete/word_0/$entry
      -- CP-element group 488: 	 branch_block_stmt_38/assign_stmt_939_to_assign_stmt_955/ptr_deref_941_Update/word_access_complete/word_0/cr
      -- CP-element group 488: 	 branch_block_stmt_38/merge_stmt_924_PhiAck/$exit
      -- CP-element group 488: 	 branch_block_stmt_38/merge_stmt_924_PhiAck/phi_stmt_925_ack
      -- 
    phi_stmt_925_ack_3649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 488_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_925_ack_0, ack => convTranspose_CP_34_elements(488)); -- 
    req_1760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(488), ack => array_obj_ref_937_index_offset_req_0); -- 
    req_1765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(488), ack => array_obj_ref_937_index_offset_req_1); -- 
    req_1780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(488), ack => addr_of_938_final_reg_req_1); -- 
    cr_1830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(488), ack => ptr_deref_941_store_0_req_1); -- 
    -- CP-element group 489:  merge  fork  transition  place  output  bypass 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	219 
    -- CP-element group 489: 	229 
    -- CP-element group 489: successors 
    -- CP-element group 489: 	231 
    -- CP-element group 489: 	232 
    -- CP-element group 489: 	234 
    -- CP-element group 489:  members (16) 
      -- CP-element group 489: 	 branch_block_stmt_38/merge_stmt_964__exit__
      -- CP-element group 489: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973__entry__
      -- CP-element group 489: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_update_start_
      -- CP-element group 489: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Sample/crr
      -- CP-element group 489: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Update/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/call_stmt_967_Update/ccr
      -- CP-element group 489: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_update_start_
      -- CP-element group 489: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Update/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/call_stmt_967_to_assign_stmt_973/type_cast_972_Update/cr
      -- CP-element group 489: 	 branch_block_stmt_38/merge_stmt_964_PhiReqMerge
      -- CP-element group 489: 	 branch_block_stmt_38/merge_stmt_964_PhiAck/$entry
      -- CP-element group 489: 	 branch_block_stmt_38/merge_stmt_964_PhiAck/$exit
      -- CP-element group 489: 	 branch_block_stmt_38/merge_stmt_964_PhiAck/dummy
      -- 
    crr_1861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(489), ack => call_stmt_967_call_req_0); -- 
    ccr_1866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(489), ack => call_stmt_967_call_req_1); -- 
    cr_1880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(489), ack => type_cast_972_inst_req_1); -- 
    convTranspose_CP_34_elements(489) <= OrReduce(convTranspose_CP_34_elements(219) & convTranspose_CP_34_elements(229));
    -- CP-element group 490:  transition  output  delay-element  bypass 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	420 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	494 
    -- CP-element group 490:  members (5) 
      -- CP-element group 490: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/$exit
      -- CP-element group 490: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1355/$exit
      -- CP-element group 490: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_sources/$exit
      -- CP-element group 490: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_sources/type_cast_1359_konst_delay_trans
      -- CP-element group 490: 	 branch_block_stmt_38/bbx_xnph_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_req
      -- 
    phi_stmt_1355_req_3695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1355_req_3695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(490), ack => phi_stmt_1355_req_0); -- 
    -- Element group convTranspose_CP_34_elements(490) is a control-delay.
    cp_element_490_delay: control_delay_element  generic map(name => " 490_delay", delay_value => 1)  port map(req => convTranspose_CP_34_elements(420), ack => convTranspose_CP_34_elements(490), clk => clk, reset =>reset);
    -- CP-element group 491:  transition  input  bypass 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	468 
    -- CP-element group 491: successors 
    -- CP-element group 491: 	493 
    -- CP-element group 491:  members (2) 
      -- CP-element group 491: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_sources/type_cast_1361/SplitProtocol/Sample/$exit
      -- CP-element group 491: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_sources/type_cast_1361/SplitProtocol/Sample/ra
      -- 
    ra_3715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 491_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1361_inst_ack_0, ack => convTranspose_CP_34_elements(491)); -- 
    -- CP-element group 492:  transition  input  bypass 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	468 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	493 
    -- CP-element group 492:  members (2) 
      -- CP-element group 492: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_sources/type_cast_1361/SplitProtocol/Update/$exit
      -- CP-element group 492: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_sources/type_cast_1361/SplitProtocol/Update/ca
      -- 
    ca_3720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1361_inst_ack_1, ack => convTranspose_CP_34_elements(492)); -- 
    -- CP-element group 493:  join  transition  output  bypass 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	491 
    -- CP-element group 493: 	492 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	494 
    -- CP-element group 493:  members (6) 
      -- CP-element group 493: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/$exit
      -- CP-element group 493: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1355/$exit
      -- CP-element group 493: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_sources/$exit
      -- CP-element group 493: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_sources/type_cast_1361/$exit
      -- CP-element group 493: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_sources/type_cast_1361/SplitProtocol/$exit
      -- CP-element group 493: 	 branch_block_stmt_38/forx_xbody427_forx_xbody427_PhiReq/phi_stmt_1355/phi_stmt_1355_req
      -- 
    phi_stmt_1355_req_3721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1355_req_3721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(493), ack => phi_stmt_1355_req_1); -- 
    convTranspose_cp_element_group_493: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_493"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_34_elements(491) & convTranspose_CP_34_elements(492);
      gj_convTranspose_cp_element_group_493 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_34_elements(493), clk => clk, reset => reset); --
    end block;
    -- CP-element group 494:  merge  transition  place  bypass 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	490 
    -- CP-element group 494: 	493 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	495 
    -- CP-element group 494:  members (2) 
      -- CP-element group 494: 	 branch_block_stmt_38/merge_stmt_1354_PhiReqMerge
      -- CP-element group 494: 	 branch_block_stmt_38/merge_stmt_1354_PhiAck/$entry
      -- 
    convTranspose_CP_34_elements(494) <= OrReduce(convTranspose_CP_34_elements(490) & convTranspose_CP_34_elements(493));
    -- CP-element group 495:  fork  transition  place  input  output  bypass 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	494 
    -- CP-element group 495: successors 
    -- CP-element group 495: 	421 
    -- CP-element group 495: 	422 
    -- CP-element group 495: 	424 
    -- CP-element group 495: 	426 
    -- CP-element group 495: 	428 
    -- CP-element group 495: 	430 
    -- CP-element group 495: 	432 
    -- CP-element group 495: 	434 
    -- CP-element group 495: 	436 
    -- CP-element group 495: 	438 
    -- CP-element group 495: 	440 
    -- CP-element group 495: 	442 
    -- CP-element group 495:  members (53) 
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1376_update_start_
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_index_resize_1/index_resize_ack
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_index_scale_1/$entry
      -- CP-element group 495: 	 branch_block_stmt_38/merge_stmt_1354__exit__
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482__entry__
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1396_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_index_scaled_1
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1396_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_final_index_sum_regn_update_start
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_index_resize_1/$entry
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_index_resized_1
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1436_update_start_
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_index_resize_1/index_resize_req
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_index_resize_1/$exit
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1426_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_index_scale_1/scale_rename_req
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1426_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/$entry
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/addr_of_1368_update_start_
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_final_index_sum_regn_Sample/$entry
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1406_update_start_
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1426_update_start_
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_index_scale_1/scale_rename_ack
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_index_computed_1
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1396_update_start_
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Update/word_access_complete/word_0/cr
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_final_index_sum_regn_Sample/req
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Update/word_access_complete/word_0/$entry
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Update/word_access_complete/$entry
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1386_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1446_update_start_
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1386_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1416_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1416_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1386_update_start_
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1376_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1416_update_start_
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/ptr_deref_1372_update_start_
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1406_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/addr_of_1368_complete/req
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1436_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/addr_of_1368_complete/$entry
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1376_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1436_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1406_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_index_scale_1/$exit
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_final_index_sum_regn_Update/req
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1446_Update/cr
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/array_obj_ref_1367_final_index_sum_regn_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_38/assign_stmt_1369_to_assign_stmt_1482/type_cast_1446_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_38/merge_stmt_1354_PhiAck/$exit
      -- CP-element group 495: 	 branch_block_stmt_38/merge_stmt_1354_PhiAck/phi_stmt_1355_ack
      -- 
    phi_stmt_1355_ack_3726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 495_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1355_ack_0, ack => convTranspose_CP_34_elements(495)); -- 
    cr_3239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(495), ack => type_cast_1396_inst_req_1); -- 
    cr_3281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(495), ack => type_cast_1426_inst_req_1); -- 
    cr_3192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(495), ack => ptr_deref_1372_load_0_req_1); -- 
    req_3127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(495), ack => array_obj_ref_1367_index_offset_req_0); -- 
    cr_3225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(495), ack => type_cast_1386_inst_req_1); -- 
    cr_3267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(495), ack => type_cast_1416_inst_req_1); -- 
    cr_3211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(495), ack => type_cast_1376_inst_req_1); -- 
    cr_3253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(495), ack => type_cast_1406_inst_req_1); -- 
    req_3147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(495), ack => addr_of_1368_final_reg_req_1); -- 
    cr_3295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(495), ack => type_cast_1436_inst_req_1); -- 
    req_3132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(495), ack => array_obj_ref_1367_index_offset_req_1); -- 
    cr_3309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_34_elements(495), ack => type_cast_1446_inst_req_1); -- 
    -- CP-element group 496:  merge  transition  place  bypass 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	418 
    -- CP-element group 496: 	467 
    -- CP-element group 496: successors 
    -- CP-element group 496:  members (16) 
      -- CP-element group 496: 	 $exit
      -- CP-element group 496: 	 branch_block_stmt_38/$exit
      -- CP-element group 496: 	 branch_block_stmt_38/branch_block_stmt_38__exit__
      -- CP-element group 496: 	 branch_block_stmt_38/merge_stmt_1491__exit__
      -- CP-element group 496: 	 branch_block_stmt_38/return__
      -- CP-element group 496: 	 branch_block_stmt_38/merge_stmt_1493__exit__
      -- CP-element group 496: 	 branch_block_stmt_38/merge_stmt_1491_PhiReqMerge
      -- CP-element group 496: 	 branch_block_stmt_38/merge_stmt_1491_PhiAck/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/merge_stmt_1491_PhiAck/$exit
      -- CP-element group 496: 	 branch_block_stmt_38/merge_stmt_1491_PhiAck/dummy
      -- CP-element group 496: 	 branch_block_stmt_38/return___PhiReq/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/return___PhiReq/$exit
      -- CP-element group 496: 	 branch_block_stmt_38/merge_stmt_1493_PhiReqMerge
      -- CP-element group 496: 	 branch_block_stmt_38/merge_stmt_1493_PhiAck/$entry
      -- CP-element group 496: 	 branch_block_stmt_38/merge_stmt_1493_PhiAck/$exit
      -- CP-element group 496: 	 branch_block_stmt_38/merge_stmt_1493_PhiAck/dummy
      -- 
    convTranspose_CP_34_elements(496) <= OrReduce(convTranspose_CP_34_elements(418) & convTranspose_CP_34_elements(467));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar525_936_resized : std_logic_vector(13 downto 0);
    signal R_indvar525_936_scaled : std_logic_vector(13 downto 0);
    signal R_indvar539_692_resized : std_logic_vector(10 downto 0);
    signal R_indvar539_692_scaled : std_logic_vector(10 downto 0);
    signal R_indvar555_485_resized : std_logic_vector(13 downto 0);
    signal R_indvar555_485_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1366_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1366_scaled : std_logic_vector(13 downto 0);
    signal add108_339 : std_logic_vector(15 downto 0);
    signal add117_364 : std_logic_vector(15 downto 0);
    signal add126_389 : std_logic_vector(15 downto 0);
    signal add12_88 : std_logic_vector(15 downto 0);
    signal add135_414 : std_logic_vector(15 downto 0);
    signal add150_513 : std_logic_vector(63 downto 0);
    signal add156_531 : std_logic_vector(63 downto 0);
    signal add162_549 : std_logic_vector(63 downto 0);
    signal add168_567 : std_logic_vector(63 downto 0);
    signal add174_585 : std_logic_vector(63 downto 0);
    signal add180_603 : std_logic_vector(63 downto 0);
    signal add186_621 : std_logic_vector(63 downto 0);
    signal add206_720 : std_logic_vector(63 downto 0);
    signal add212_738 : std_logic_vector(63 downto 0);
    signal add218_756 : std_logic_vector(63 downto 0);
    signal add21_113 : std_logic_vector(15 downto 0);
    signal add224_774 : std_logic_vector(63 downto 0);
    signal add230_792 : std_logic_vector(63 downto 0);
    signal add236_810 : std_logic_vector(63 downto 0);
    signal add242_828 : std_logic_vector(63 downto 0);
    signal add30_138 : std_logic_vector(15 downto 0);
    signal add39_163 : std_logic_vector(15 downto 0);
    signal add48_188 : std_logic_vector(15 downto 0);
    signal add57_213 : std_logic_vector(15 downto 0);
    signal add74_253 : std_logic_vector(31 downto 0);
    signal add79_258 : std_logic_vector(31 downto 0);
    signal add99_314 : std_logic_vector(15 downto 0);
    signal add_63 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1367_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1367_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1367_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1367_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1367_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1367_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_486_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_486_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_486_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_486_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_486_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_486_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_693_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_693_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_693_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_693_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_693_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_693_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_937_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_937_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_937_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_937_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_937_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_937_root_address : std_logic_vector(13 downto 0);
    signal arrayidx246_695 : std_logic_vector(31 downto 0);
    signal arrayidx269_939 : std_logic_vector(31 downto 0);
    signal arrayidx432_1369 : std_logic_vector(31 downto 0);
    signal arrayidx_488 : std_logic_vector(31 downto 0);
    signal call101_317 : std_logic_vector(7 downto 0);
    signal call106_330 : std_logic_vector(7 downto 0);
    signal call10_79 : std_logic_vector(7 downto 0);
    signal call110_342 : std_logic_vector(7 downto 0);
    signal call115_355 : std_logic_vector(7 downto 0);
    signal call119_367 : std_logic_vector(7 downto 0);
    signal call124_380 : std_logic_vector(7 downto 0);
    signal call128_392 : std_logic_vector(7 downto 0);
    signal call133_405 : std_logic_vector(7 downto 0);
    signal call143_491 : std_logic_vector(7 downto 0);
    signal call147_504 : std_logic_vector(7 downto 0);
    signal call14_91 : std_logic_vector(7 downto 0);
    signal call153_522 : std_logic_vector(7 downto 0);
    signal call159_540 : std_logic_vector(7 downto 0);
    signal call165_558 : std_logic_vector(7 downto 0);
    signal call171_576 : std_logic_vector(7 downto 0);
    signal call177_594 : std_logic_vector(7 downto 0);
    signal call183_612 : std_logic_vector(7 downto 0);
    signal call199_698 : std_logic_vector(7 downto 0);
    signal call19_104 : std_logic_vector(7 downto 0);
    signal call203_711 : std_logic_vector(7 downto 0);
    signal call209_729 : std_logic_vector(7 downto 0);
    signal call215_747 : std_logic_vector(7 downto 0);
    signal call221_765 : std_logic_vector(7 downto 0);
    signal call227_783 : std_logic_vector(7 downto 0);
    signal call233_801 : std_logic_vector(7 downto 0);
    signal call239_819 : std_logic_vector(7 downto 0);
    signal call23_116 : std_logic_vector(7 downto 0);
    signal call275_967 : std_logic_vector(63 downto 0);
    signal call28_129 : std_logic_vector(7 downto 0);
    signal call2_54 : std_logic_vector(7 downto 0);
    signal call32_141 : std_logic_vector(7 downto 0);
    signal call346_1189 : std_logic_vector(15 downto 0);
    signal call348_1192 : std_logic_vector(15 downto 0);
    signal call350_1195 : std_logic_vector(15 downto 0);
    signal call352_1198 : std_logic_vector(15 downto 0);
    signal call354_1201 : std_logic_vector(63 downto 0);
    signal call37_154 : std_logic_vector(7 downto 0);
    signal call41_166 : std_logic_vector(7 downto 0);
    signal call46_179 : std_logic_vector(7 downto 0);
    signal call50_191 : std_logic_vector(7 downto 0);
    signal call55_204 : std_logic_vector(7 downto 0);
    signal call5_66 : std_logic_vector(7 downto 0);
    signal call92_292 : std_logic_vector(7 downto 0);
    signal call97_305 : std_logic_vector(7 downto 0);
    signal call_41 : std_logic_vector(7 downto 0);
    signal cmp194509_435 : std_logic_vector(0 downto 0);
    signal cmp264505_880 : std_logic_vector(0 downto 0);
    signal cmp513_420 : std_logic_vector(0 downto 0);
    signal conv104_321 : std_logic_vector(15 downto 0);
    signal conv107_334 : std_logic_vector(15 downto 0);
    signal conv113_346 : std_logic_vector(15 downto 0);
    signal conv116_359 : std_logic_vector(15 downto 0);
    signal conv11_83 : std_logic_vector(15 downto 0);
    signal conv122_371 : std_logic_vector(15 downto 0);
    signal conv125_384 : std_logic_vector(15 downto 0);
    signal conv131_396 : std_logic_vector(15 downto 0);
    signal conv134_409 : std_logic_vector(15 downto 0);
    signal conv144_495 : std_logic_vector(63 downto 0);
    signal conv149_508 : std_logic_vector(63 downto 0);
    signal conv155_526 : std_logic_vector(63 downto 0);
    signal conv161_544 : std_logic_vector(63 downto 0);
    signal conv167_562 : std_logic_vector(63 downto 0);
    signal conv173_580 : std_logic_vector(63 downto 0);
    signal conv179_598 : std_logic_vector(63 downto 0);
    signal conv17_95 : std_logic_vector(15 downto 0);
    signal conv185_616 : std_logic_vector(63 downto 0);
    signal conv1_45 : std_logic_vector(15 downto 0);
    signal conv200_702 : std_logic_vector(63 downto 0);
    signal conv205_715 : std_logic_vector(63 downto 0);
    signal conv20_108 : std_logic_vector(15 downto 0);
    signal conv211_733 : std_logic_vector(63 downto 0);
    signal conv217_751 : std_logic_vector(63 downto 0);
    signal conv223_769 : std_logic_vector(63 downto 0);
    signal conv229_787 : std_logic_vector(63 downto 0);
    signal conv235_805 : std_logic_vector(63 downto 0);
    signal conv241_823 : std_logic_vector(63 downto 0);
    signal conv253_856 : std_logic_vector(31 downto 0);
    signal conv255_860 : std_logic_vector(31 downto 0);
    signal conv258_864 : std_logic_vector(31 downto 0);
    signal conv26_120 : std_logic_vector(15 downto 0);
    signal conv276_973 : std_logic_vector(63 downto 0);
    signal conv29_133 : std_logic_vector(15 downto 0);
    signal conv305_1055 : std_logic_vector(15 downto 0);
    signal conv307_1062 : std_logic_vector(15 downto 0);
    signal conv322_1111 : std_logic_vector(15 downto 0);
    signal conv324_1118 : std_logic_vector(15 downto 0);
    signal conv339_1167 : std_logic_vector(15 downto 0);
    signal conv341_1174 : std_logic_vector(15 downto 0);
    signal conv355_1206 : std_logic_vector(63 downto 0);
    signal conv35_145 : std_logic_vector(15 downto 0);
    signal conv361_1215 : std_logic_vector(7 downto 0);
    signal conv367_1225 : std_logic_vector(7 downto 0);
    signal conv373_1235 : std_logic_vector(7 downto 0);
    signal conv379_1245 : std_logic_vector(7 downto 0);
    signal conv385_1255 : std_logic_vector(7 downto 0);
    signal conv38_158 : std_logic_vector(15 downto 0);
    signal conv391_1265 : std_logic_vector(7 downto 0);
    signal conv397_1275 : std_logic_vector(7 downto 0);
    signal conv3_58 : std_logic_vector(15 downto 0);
    signal conv403_1285 : std_logic_vector(7 downto 0);
    signal conv437_1377 : std_logic_vector(7 downto 0);
    signal conv443_1387 : std_logic_vector(7 downto 0);
    signal conv449_1397 : std_logic_vector(7 downto 0);
    signal conv44_170 : std_logic_vector(15 downto 0);
    signal conv455_1407 : std_logic_vector(7 downto 0);
    signal conv461_1417 : std_logic_vector(7 downto 0);
    signal conv467_1427 : std_logic_vector(7 downto 0);
    signal conv473_1437 : std_logic_vector(7 downto 0);
    signal conv479_1447 : std_logic_vector(7 downto 0);
    signal conv47_183 : std_logic_vector(15 downto 0);
    signal conv53_195 : std_logic_vector(15 downto 0);
    signal conv56_208 : std_logic_vector(15 downto 0);
    signal conv61_217 : std_logic_vector(31 downto 0);
    signal conv63_221 : std_logic_vector(31 downto 0);
    signal conv65_225 : std_logic_vector(31 downto 0);
    signal conv82_262 : std_logic_vector(31 downto 0);
    signal conv84_266 : std_logic_vector(31 downto 0);
    signal conv87_270 : std_logic_vector(31 downto 0);
    signal conv8_70 : std_logic_vector(15 downto 0);
    signal conv90_274 : std_logic_vector(31 downto 0);
    signal conv95_296 : std_logic_vector(15 downto 0);
    signal conv98_309 : std_logic_vector(15 downto 0);
    signal exitcond1_1482 : std_logic_vector(0 downto 0);
    signal exitcond2_843 : std_logic_vector(0 downto 0);
    signal exitcond3_636 : std_logic_vector(0 downto 0);
    signal exitcond_955 : std_logic_vector(0 downto 0);
    signal iNsTr_14_247 : std_logic_vector(31 downto 0);
    signal iNsTr_195_1339 : std_logic_vector(63 downto 0);
    signal iNsTr_26_458 : std_logic_vector(63 downto 0);
    signal iNsTr_39_665 : std_logic_vector(63 downto 0);
    signal iNsTr_53_909 : std_logic_vector(63 downto 0);
    signal indvar525_925 : std_logic_vector(63 downto 0);
    signal indvar539_681 : std_logic_vector(63 downto 0);
    signal indvar555_474 : std_logic_vector(63 downto 0);
    signal indvar_1355 : std_logic_vector(63 downto 0);
    signal indvarx_xnext526_950 : std_logic_vector(63 downto 0);
    signal indvarx_xnext540_838 : std_logic_vector(63 downto 0);
    signal indvarx_xnext556_631 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1477 : std_logic_vector(63 downto 0);
    signal mul256_869 : std_logic_vector(31 downto 0);
    signal mul259_874 : std_logic_vector(31 downto 0);
    signal mul66_235 : std_logic_vector(31 downto 0);
    signal mul85_279 : std_logic_vector(31 downto 0);
    signal mul88_284 : std_logic_vector(31 downto 0);
    signal mul91_289 : std_logic_vector(31 downto 0);
    signal mul_230 : std_logic_vector(31 downto 0);
    signal ptr_deref_1372_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1372_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1372_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1372_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1372_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_623_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_623_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_623_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_623_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_623_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_623_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_830_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_830_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_830_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_830_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_830_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_830_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_941_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_941_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_941_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_941_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_941_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_941_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl105_327 : std_logic_vector(15 downto 0);
    signal shl114_352 : std_logic_vector(15 downto 0);
    signal shl123_377 : std_logic_vector(15 downto 0);
    signal shl132_402 : std_logic_vector(15 downto 0);
    signal shl146_501 : std_logic_vector(63 downto 0);
    signal shl152_519 : std_logic_vector(63 downto 0);
    signal shl158_537 : std_logic_vector(63 downto 0);
    signal shl164_555 : std_logic_vector(63 downto 0);
    signal shl170_573 : std_logic_vector(63 downto 0);
    signal shl176_591 : std_logic_vector(63 downto 0);
    signal shl182_609 : std_logic_vector(63 downto 0);
    signal shl18_101 : std_logic_vector(15 downto 0);
    signal shl202_708 : std_logic_vector(63 downto 0);
    signal shl208_726 : std_logic_vector(63 downto 0);
    signal shl214_744 : std_logic_vector(63 downto 0);
    signal shl220_762 : std_logic_vector(63 downto 0);
    signal shl226_780 : std_logic_vector(63 downto 0);
    signal shl232_798 : std_logic_vector(63 downto 0);
    signal shl238_816 : std_logic_vector(63 downto 0);
    signal shl27_126 : std_logic_vector(15 downto 0);
    signal shl36_151 : std_logic_vector(15 downto 0);
    signal shl45_176 : std_logic_vector(15 downto 0);
    signal shl54_201 : std_logic_vector(15 downto 0);
    signal shl96_302 : std_logic_vector(15 downto 0);
    signal shl9_76 : std_logic_vector(15 downto 0);
    signal shl_51 : std_logic_vector(15 downto 0);
    signal shr304_1051 : std_logic_vector(31 downto 0);
    signal shr321_1107 : std_logic_vector(31 downto 0);
    signal shr338_1163 : std_logic_vector(31 downto 0);
    signal shr364_1221 : std_logic_vector(63 downto 0);
    signal shr370_1231 : std_logic_vector(63 downto 0);
    signal shr376_1241 : std_logic_vector(63 downto 0);
    signal shr382_1251 : std_logic_vector(63 downto 0);
    signal shr388_1261 : std_logic_vector(63 downto 0);
    signal shr394_1271 : std_logic_vector(63 downto 0);
    signal shr400_1281 : std_logic_vector(63 downto 0);
    signal shr440_1383 : std_logic_vector(63 downto 0);
    signal shr446_1393 : std_logic_vector(63 downto 0);
    signal shr452_1403 : std_logic_vector(63 downto 0);
    signal shr458_1413 : std_logic_vector(63 downto 0);
    signal shr464_1423 : std_logic_vector(63 downto 0);
    signal shr470_1433 : std_logic_vector(63 downto 0);
    signal shr476_1443 : std_logic_vector(63 downto 0);
    signal shr_241 : std_logic_vector(31 downto 0);
    signal sub_1211 : std_logic_vector(63 downto 0);
    signal tmp433_1373 : std_logic_vector(63 downto 0);
    signal tmp520_1323 : std_logic_vector(31 downto 0);
    signal tmp520x_xop_1335 : std_logic_vector(31 downto 0);
    signal tmp521_1329 : std_logic_vector(0 downto 0);
    signal tmp524_1352 : std_logic_vector(63 downto 0);
    signal tmp532_893 : std_logic_vector(31 downto 0);
    signal tmp532x_xop_905 : std_logic_vector(31 downto 0);
    signal tmp533_899 : std_logic_vector(0 downto 0);
    signal tmp537_922 : std_logic_vector(63 downto 0);
    signal tmp548_649 : std_logic_vector(31 downto 0);
    signal tmp548x_xop_661 : std_logic_vector(31 downto 0);
    signal tmp549_655 : std_logic_vector(0 downto 0);
    signal tmp553_678 : std_logic_vector(63 downto 0);
    signal tmp562x_xop_454 : std_logic_vector(31 downto 0);
    signal tmp563_448 : std_logic_vector(0 downto 0);
    signal tmp567_471 : std_logic_vector(63 downto 0);
    signal type_cast_1004_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1008_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1049_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1105_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1161_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1204_wire : std_logic_vector(63 downto 0);
    signal type_cast_1219_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1229_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1239_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1249_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_124_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1259_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1269_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1279_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1321_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1327_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1333_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1343_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1350_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1359_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1361_wire : std_logic_vector(63 downto 0);
    signal type_cast_1381_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1391_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1401_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1411_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1421_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1431_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1441_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1475_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_149_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_174_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_199_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_239_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_245_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_251_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_300_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_325_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_350_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_375_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_400_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_418_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_433_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_446_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_452_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_462_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_469_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_478_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_480_wire : std_logic_vector(63 downto 0);
    signal type_cast_499_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_49_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_517_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_535_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_553_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_571_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_589_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_607_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_629_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_647_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_653_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_659_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_669_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_676_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_685_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_687_wire : std_logic_vector(63 downto 0);
    signal type_cast_706_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_724_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_742_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_74_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_760_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_778_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_796_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_814_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_836_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_878_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_891_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_897_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_903_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_913_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_920_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_928_wire : std_logic_vector(63 downto 0);
    signal type_cast_931_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_943_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_948_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_971_wire : std_logic_vector(63 downto 0);
    signal type_cast_99_wire_constant : std_logic_vector(15 downto 0);
    signal xx_xop569_915 : std_logic_vector(63 downto 0);
    signal xx_xop570_671 : std_logic_vector(63 downto 0);
    signal xx_xop571_464 : std_logic_vector(63 downto 0);
    signal xx_xop_1345 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1367_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1367_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1367_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1367_resized_base_address <= "00000000000000";
    array_obj_ref_486_constant_part_of_offset <= "00000000000000";
    array_obj_ref_486_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_486_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_486_resized_base_address <= "00000000000000";
    array_obj_ref_693_constant_part_of_offset <= "00000100010";
    array_obj_ref_693_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_693_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_693_resized_base_address <= "00000000000";
    array_obj_ref_937_constant_part_of_offset <= "00000000000000";
    array_obj_ref_937_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_937_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_937_resized_base_address <= "00000000000000";
    ptr_deref_1372_word_offset_0 <= "00000000000000";
    ptr_deref_623_word_offset_0 <= "00000000000000";
    ptr_deref_830_word_offset_0 <= "00000000000";
    ptr_deref_941_word_offset_0 <= "00000000000000";
    type_cast_1004_wire_constant <= "0000000000000000";
    type_cast_1008_wire_constant <= "0000000000000000";
    type_cast_1049_wire_constant <= "00000000000000000000000000010010";
    type_cast_1105_wire_constant <= "00000000000000000000000000010001";
    type_cast_1161_wire_constant <= "00000000000000000000000000010000";
    type_cast_1219_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1229_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1239_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1249_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_124_wire_constant <= "0000000000001000";
    type_cast_1259_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1269_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1279_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1321_wire_constant <= "00000000000000000000000000000010";
    type_cast_1327_wire_constant <= "00000000000000000000000000000001";
    type_cast_1333_wire_constant <= "11111111111111111111111111111111";
    type_cast_1343_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1350_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1359_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1381_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1391_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1401_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1411_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1421_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1431_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1441_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1475_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_149_wire_constant <= "0000000000001000";
    type_cast_174_wire_constant <= "0000000000001000";
    type_cast_199_wire_constant <= "0000000000001000";
    type_cast_239_wire_constant <= "00000000000000000000000000000010";
    type_cast_245_wire_constant <= "00000000000000000000000000000001";
    type_cast_251_wire_constant <= "01111111111111111111111111111110";
    type_cast_300_wire_constant <= "0000000000001000";
    type_cast_325_wire_constant <= "0000000000001000";
    type_cast_350_wire_constant <= "0000000000001000";
    type_cast_375_wire_constant <= "0000000000001000";
    type_cast_400_wire_constant <= "0000000000001000";
    type_cast_418_wire_constant <= "00000000000000000000000000000011";
    type_cast_433_wire_constant <= "00000000000000000000000000000011";
    type_cast_446_wire_constant <= "00000000000000000000000000000001";
    type_cast_452_wire_constant <= "11111111111111111111111111111111";
    type_cast_462_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_469_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_478_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_499_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_49_wire_constant <= "0000000000001000";
    type_cast_517_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_535_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_553_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_571_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_589_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_607_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_629_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_647_wire_constant <= "00000000000000000000000000000010";
    type_cast_653_wire_constant <= "00000000000000000000000000000001";
    type_cast_659_wire_constant <= "11111111111111111111111111111111";
    type_cast_669_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_676_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_685_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_706_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_724_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_742_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_74_wire_constant <= "0000000000001000";
    type_cast_760_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_778_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_796_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_814_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_836_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_878_wire_constant <= "00000000000000000000000000000011";
    type_cast_891_wire_constant <= "00000000000000000000000000000010";
    type_cast_897_wire_constant <= "00000000000000000000000000000001";
    type_cast_903_wire_constant <= "11111111111111111111111111111111";
    type_cast_913_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_920_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_931_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_943_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_948_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_99_wire_constant <= "0000000000001000";
    phi_stmt_1355: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1359_wire_constant & type_cast_1361_wire;
      req <= phi_stmt_1355_req_0 & phi_stmt_1355_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1355",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1355_ack_0,
          idata => idata,
          odata => indvar_1355,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1355
    phi_stmt_474: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_478_wire_constant & type_cast_480_wire;
      req <= phi_stmt_474_req_0 & phi_stmt_474_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_474",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_474_ack_0,
          idata => idata,
          odata => indvar555_474,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_474
    phi_stmt_681: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_685_wire_constant & type_cast_687_wire;
      req <= phi_stmt_681_req_0 & phi_stmt_681_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_681",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_681_ack_0,
          idata => idata,
          odata => indvar539_681,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_681
    phi_stmt_925: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_928_wire & type_cast_931_wire_constant;
      req <= phi_stmt_925_req_0 & phi_stmt_925_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_925",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_925_ack_0,
          idata => idata,
          odata => indvar525_925,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_925
    -- flow-through select operator MUX_1351_inst
    tmp524_1352 <= xx_xop_1345 when (tmp521_1329(0) /=  '0') else type_cast_1350_wire_constant;
    -- flow-through select operator MUX_470_inst
    tmp567_471 <= xx_xop571_464 when (tmp563_448(0) /=  '0') else type_cast_469_wire_constant;
    -- flow-through select operator MUX_677_inst
    tmp553_678 <= xx_xop570_671 when (tmp549_655(0) /=  '0') else type_cast_676_wire_constant;
    -- flow-through select operator MUX_921_inst
    tmp537_922 <= xx_xop569_915 when (tmp533_899(0) /=  '0') else type_cast_920_wire_constant;
    addr_of_1368_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1368_final_reg_req_0;
      addr_of_1368_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1368_final_reg_req_1;
      addr_of_1368_final_reg_ack_1<= rack(0);
      addr_of_1368_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1368_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1367_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx432_1369,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_487_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_487_final_reg_req_0;
      addr_of_487_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_487_final_reg_req_1;
      addr_of_487_final_reg_ack_1<= rack(0);
      addr_of_487_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_487_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_486_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_488,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_694_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_694_final_reg_req_0;
      addr_of_694_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_694_final_reg_req_1;
      addr_of_694_final_reg_ack_1<= rack(0);
      addr_of_694_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_694_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_693_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx246_695,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_938_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_938_final_reg_req_0;
      addr_of_938_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_938_final_reg_req_1;
      addr_of_938_final_reg_ack_1<= rack(0);
      addr_of_938_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_938_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_937_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx269_939,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1054_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1054_inst_req_0;
      type_cast_1054_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1054_inst_req_1;
      type_cast_1054_inst_ack_1<= rack(0);
      type_cast_1054_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1054_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr304_1051,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv305_1055,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1061_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1061_inst_req_0;
      type_cast_1061_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1061_inst_req_1;
      type_cast_1061_inst_ack_1<= rack(0);
      type_cast_1061_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1061_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_241,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv307_1062,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_107_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_107_inst_req_0;
      type_cast_107_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_107_inst_req_1;
      type_cast_107_inst_ack_1<= rack(0);
      type_cast_107_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_107_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_104,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_108,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1110_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1110_inst_req_0;
      type_cast_1110_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1110_inst_req_1;
      type_cast_1110_inst_ack_1<= rack(0);
      type_cast_1110_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1110_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr321_1107,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv322_1111,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1117_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1117_inst_req_0;
      type_cast_1117_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1117_inst_req_1;
      type_cast_1117_inst_ack_1<= rack(0);
      type_cast_1117_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1117_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add74_253,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv324_1118,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1166_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1166_inst_req_0;
      type_cast_1166_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1166_inst_req_1;
      type_cast_1166_inst_ack_1<= rack(0);
      type_cast_1166_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1166_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr338_1163,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv339_1167,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1173_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1173_inst_req_0;
      type_cast_1173_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1173_inst_req_1;
      type_cast_1173_inst_ack_1<= rack(0);
      type_cast_1173_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1173_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add79_258,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv341_1174,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_119_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_119_inst_req_0;
      type_cast_119_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_119_inst_req_1;
      type_cast_119_inst_ack_1<= rack(0);
      type_cast_119_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_119_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_116,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_120,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1205_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1205_inst_req_0;
      type_cast_1205_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1205_inst_req_1;
      type_cast_1205_inst_ack_1<= rack(0);
      type_cast_1205_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1205_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1204_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv355_1206,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1214_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1214_inst_req_0;
      type_cast_1214_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1214_inst_req_1;
      type_cast_1214_inst_ack_1<= rack(0);
      type_cast_1214_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1214_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1211,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv361_1215,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1224_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1224_inst_req_0;
      type_cast_1224_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1224_inst_req_1;
      type_cast_1224_inst_ack_1<= rack(0);
      type_cast_1224_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1224_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr364_1221,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv367_1225,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1234_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1234_inst_req_0;
      type_cast_1234_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1234_inst_req_1;
      type_cast_1234_inst_ack_1<= rack(0);
      type_cast_1234_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1234_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr370_1231,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv373_1235,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1244_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1244_inst_req_0;
      type_cast_1244_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1244_inst_req_1;
      type_cast_1244_inst_ack_1<= rack(0);
      type_cast_1244_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1244_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr376_1241,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv379_1245,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1254_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1254_inst_req_0;
      type_cast_1254_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1254_inst_req_1;
      type_cast_1254_inst_ack_1<= rack(0);
      type_cast_1254_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1254_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr382_1251,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv385_1255,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1264_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1264_inst_req_0;
      type_cast_1264_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1264_inst_req_1;
      type_cast_1264_inst_ack_1<= rack(0);
      type_cast_1264_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1264_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr388_1261,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv391_1265,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1274_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1274_inst_req_0;
      type_cast_1274_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1274_inst_req_1;
      type_cast_1274_inst_ack_1<= rack(0);
      type_cast_1274_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1274_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr394_1271,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv397_1275,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1284_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1284_inst_req_0;
      type_cast_1284_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1284_inst_req_1;
      type_cast_1284_inst_ack_1<= rack(0);
      type_cast_1284_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1284_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr400_1281,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv403_1285,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_132_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_132_inst_req_0;
      type_cast_132_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_132_inst_req_1;
      type_cast_132_inst_ack_1<= rack(0);
      type_cast_132_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_132_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_129,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_133,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1338_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1338_inst_req_0;
      type_cast_1338_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1338_inst_req_1;
      type_cast_1338_inst_ack_1<= rack(0);
      type_cast_1338_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1338_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp520x_xop_1335,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_195_1339,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1361_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1361_inst_req_0;
      type_cast_1361_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1361_inst_req_1;
      type_cast_1361_inst_ack_1<= rack(0);
      type_cast_1361_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1361_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1477,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1361_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1376_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1376_inst_req_0;
      type_cast_1376_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1376_inst_req_1;
      type_cast_1376_inst_ack_1<= rack(0);
      type_cast_1376_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1376_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp433_1373,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv437_1377,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1386_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1386_inst_req_0;
      type_cast_1386_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1386_inst_req_1;
      type_cast_1386_inst_ack_1<= rack(0);
      type_cast_1386_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1386_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr440_1383,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv443_1387,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1396_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1396_inst_req_0;
      type_cast_1396_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1396_inst_req_1;
      type_cast_1396_inst_ack_1<= rack(0);
      type_cast_1396_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1396_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr446_1393,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv449_1397,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1406_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1406_inst_req_0;
      type_cast_1406_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1406_inst_req_1;
      type_cast_1406_inst_ack_1<= rack(0);
      type_cast_1406_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1406_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr452_1403,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv455_1407,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1416_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1416_inst_req_0;
      type_cast_1416_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1416_inst_req_1;
      type_cast_1416_inst_ack_1<= rack(0);
      type_cast_1416_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1416_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr458_1413,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv461_1417,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1426_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1426_inst_req_0;
      type_cast_1426_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1426_inst_req_1;
      type_cast_1426_inst_ack_1<= rack(0);
      type_cast_1426_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1426_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr464_1423,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv467_1427,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1436_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1436_inst_req_0;
      type_cast_1436_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1436_inst_req_1;
      type_cast_1436_inst_ack_1<= rack(0);
      type_cast_1436_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1436_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr470_1433,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv473_1437,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1446_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1446_inst_req_0;
      type_cast_1446_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1446_inst_req_1;
      type_cast_1446_inst_ack_1<= rack(0);
      type_cast_1446_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1446_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr476_1443,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv479_1447,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_144_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_144_inst_req_0;
      type_cast_144_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_144_inst_req_1;
      type_cast_144_inst_ack_1<= rack(0);
      type_cast_144_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_144_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_141,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_145,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_157_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_157_inst_req_0;
      type_cast_157_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_157_inst_req_1;
      type_cast_157_inst_ack_1<= rack(0);
      type_cast_157_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_157_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_154,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_158,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_169_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_169_inst_req_0;
      type_cast_169_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_169_inst_req_1;
      type_cast_169_inst_ack_1<= rack(0);
      type_cast_169_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_169_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_166,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_170,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_182_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_182_inst_req_0;
      type_cast_182_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_182_inst_req_1;
      type_cast_182_inst_ack_1<= rack(0);
      type_cast_182_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_182_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_179,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_183,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_194_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_194_inst_req_0;
      type_cast_194_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_194_inst_req_1;
      type_cast_194_inst_ack_1<= rack(0);
      type_cast_194_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_194_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_191,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_195,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_207_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_207_inst_req_0;
      type_cast_207_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_207_inst_req_1;
      type_cast_207_inst_ack_1<= rack(0);
      type_cast_207_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_207_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_204,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_208,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_216_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_216_inst_req_0;
      type_cast_216_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_216_inst_req_1;
      type_cast_216_inst_ack_1<= rack(0);
      type_cast_216_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_216_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_63,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_217,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_220_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_220_inst_req_0;
      type_cast_220_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_220_inst_req_1;
      type_cast_220_inst_ack_1<= rack(0);
      type_cast_220_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_220_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add12_88,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_221,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_224_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_224_inst_req_0;
      type_cast_224_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_224_inst_req_1;
      type_cast_224_inst_ack_1<= rack(0);
      type_cast_224_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_224_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_113,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_225,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_261_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_261_inst_req_0;
      type_cast_261_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_261_inst_req_1;
      type_cast_261_inst_ack_1<= rack(0);
      type_cast_261_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_261_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_138,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv82_262,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_265_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_265_inst_req_0;
      type_cast_265_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_265_inst_req_1;
      type_cast_265_inst_ack_1<= rack(0);
      type_cast_265_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_265_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_163,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_266,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_269_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_269_inst_req_0;
      type_cast_269_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_269_inst_req_1;
      type_cast_269_inst_ack_1<= rack(0);
      type_cast_269_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_269_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv87_270,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_273_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_273_inst_req_0;
      type_cast_273_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_273_inst_req_1;
      type_cast_273_inst_ack_1<= rack(0);
      type_cast_273_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_273_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add57_213,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_274,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_295_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_295_inst_req_0;
      type_cast_295_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_295_inst_req_1;
      type_cast_295_inst_ack_1<= rack(0);
      type_cast_295_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_295_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call92_292,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_296,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_308_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_308_inst_req_0;
      type_cast_308_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_308_inst_req_1;
      type_cast_308_inst_ack_1<= rack(0);
      type_cast_308_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_308_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_305,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_309,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_320_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_320_inst_req_0;
      type_cast_320_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_320_inst_req_1;
      type_cast_320_inst_ack_1<= rack(0);
      type_cast_320_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_320_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_317,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_321,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_333_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_333_inst_req_0;
      type_cast_333_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_333_inst_req_1;
      type_cast_333_inst_ack_1<= rack(0);
      type_cast_333_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_333_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_330,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_334,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_345_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_345_inst_req_0;
      type_cast_345_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_345_inst_req_1;
      type_cast_345_inst_ack_1<= rack(0);
      type_cast_345_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_345_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call110_342,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_346,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_358_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_358_inst_req_0;
      type_cast_358_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_358_inst_req_1;
      type_cast_358_inst_ack_1<= rack(0);
      type_cast_358_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_358_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_359,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_370_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_370_inst_req_0;
      type_cast_370_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_370_inst_req_1;
      type_cast_370_inst_ack_1<= rack(0);
      type_cast_370_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_370_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_367,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_371,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_383_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_383_inst_req_0;
      type_cast_383_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_383_inst_req_1;
      type_cast_383_inst_ack_1<= rack(0);
      type_cast_383_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_383_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_380,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_384,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_395_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_395_inst_req_0;
      type_cast_395_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_395_inst_req_1;
      type_cast_395_inst_ack_1<= rack(0);
      type_cast_395_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_395_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_396,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_408_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_408_inst_req_0;
      type_cast_408_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_408_inst_req_1;
      type_cast_408_inst_ack_1<= rack(0);
      type_cast_408_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_408_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_405,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_409,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_44_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_44_inst_req_0;
      type_cast_44_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_44_inst_req_1;
      type_cast_44_inst_ack_1<= rack(0);
      type_cast_44_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_44_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_41,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_45,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_457_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_457_inst_req_0;
      type_cast_457_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_457_inst_req_1;
      type_cast_457_inst_ack_1<= rack(0);
      type_cast_457_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_457_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp562x_xop_454,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_26_458,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_480_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_480_inst_req_0;
      type_cast_480_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_480_inst_req_1;
      type_cast_480_inst_ack_1<= rack(0);
      type_cast_480_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_480_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext556_631,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_480_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_494_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_494_inst_req_0;
      type_cast_494_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_494_inst_req_1;
      type_cast_494_inst_ack_1<= rack(0);
      type_cast_494_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_494_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call143_491,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_495,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_507_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_507_inst_req_0;
      type_cast_507_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_507_inst_req_1;
      type_cast_507_inst_ack_1<= rack(0);
      type_cast_507_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_507_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call147_504,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv149_508,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_525_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_525_inst_req_0;
      type_cast_525_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_525_inst_req_1;
      type_cast_525_inst_ack_1<= rack(0);
      type_cast_525_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_525_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call153_522,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_526,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_543_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_543_inst_req_0;
      type_cast_543_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_543_inst_req_1;
      type_cast_543_inst_ack_1<= rack(0);
      type_cast_543_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_543_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call159_540,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_544,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_561_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_561_inst_req_0;
      type_cast_561_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_561_inst_req_1;
      type_cast_561_inst_ack_1<= rack(0);
      type_cast_561_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_561_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call165_558,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv167_562,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_579_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_579_inst_req_0;
      type_cast_579_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_579_inst_req_1;
      type_cast_579_inst_ack_1<= rack(0);
      type_cast_579_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_579_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call171_576,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_580,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_57_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_57_inst_req_0;
      type_cast_57_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_57_inst_req_1;
      type_cast_57_inst_ack_1<= rack(0);
      type_cast_57_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_57_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_54,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_58,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_597_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_597_inst_req_0;
      type_cast_597_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_597_inst_req_1;
      type_cast_597_inst_ack_1<= rack(0);
      type_cast_597_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_597_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call177_594,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv179_598,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_615_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_615_inst_req_0;
      type_cast_615_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_615_inst_req_1;
      type_cast_615_inst_ack_1<= rack(0);
      type_cast_615_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_615_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call183_612,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv185_616,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_664_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_664_inst_req_0;
      type_cast_664_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_664_inst_req_1;
      type_cast_664_inst_ack_1<= rack(0);
      type_cast_664_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_664_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp548x_xop_661,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_39_665,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_687_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_687_inst_req_0;
      type_cast_687_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_687_inst_req_1;
      type_cast_687_inst_ack_1<= rack(0);
      type_cast_687_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_687_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext540_838,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_687_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_69_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_69_inst_req_0;
      type_cast_69_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_69_inst_req_1;
      type_cast_69_inst_ack_1<= rack(0);
      type_cast_69_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_69_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_66,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_70,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_701_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_701_inst_req_0;
      type_cast_701_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_701_inst_req_1;
      type_cast_701_inst_ack_1<= rack(0);
      type_cast_701_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_701_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call199_698,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_702,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_714_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_714_inst_req_0;
      type_cast_714_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_714_inst_req_1;
      type_cast_714_inst_ack_1<= rack(0);
      type_cast_714_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_714_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call203_711,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv205_715,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_732_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_732_inst_req_0;
      type_cast_732_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_732_inst_req_1;
      type_cast_732_inst_ack_1<= rack(0);
      type_cast_732_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_732_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call209_729,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv211_733,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_750_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_750_inst_req_0;
      type_cast_750_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_750_inst_req_1;
      type_cast_750_inst_ack_1<= rack(0);
      type_cast_750_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_750_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call215_747,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv217_751,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_768_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_768_inst_req_0;
      type_cast_768_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_768_inst_req_1;
      type_cast_768_inst_ack_1<= rack(0);
      type_cast_768_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_768_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call221_765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv223_769,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_786_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_786_inst_req_0;
      type_cast_786_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_786_inst_req_1;
      type_cast_786_inst_ack_1<= rack(0);
      type_cast_786_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_786_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call227_783,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv229_787,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_804_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_804_inst_req_0;
      type_cast_804_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_804_inst_req_1;
      type_cast_804_inst_ack_1<= rack(0);
      type_cast_804_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_804_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call233_801,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv235_805,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_822_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_822_inst_req_0;
      type_cast_822_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_822_inst_req_1;
      type_cast_822_inst_ack_1<= rack(0);
      type_cast_822_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_822_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call239_819,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_823,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_82_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_82_inst_req_0;
      type_cast_82_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_82_inst_req_1;
      type_cast_82_inst_ack_1<= rack(0);
      type_cast_82_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_82_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_79,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_83,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_855_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_855_inst_req_0;
      type_cast_855_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_855_inst_req_1;
      type_cast_855_inst_ack_1<= rack(0);
      type_cast_855_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_855_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add117_364,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv253_856,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_859_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_859_inst_req_0;
      type_cast_859_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_859_inst_req_1;
      type_cast_859_inst_ack_1<= rack(0);
      type_cast_859_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_859_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add126_389,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_860,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_863_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_863_inst_req_0;
      type_cast_863_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_863_inst_req_1;
      type_cast_863_inst_ack_1<= rack(0);
      type_cast_863_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_863_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add135_414,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv258_864,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_908_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_908_inst_req_0;
      type_cast_908_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_908_inst_req_1;
      type_cast_908_inst_ack_1<= rack(0);
      type_cast_908_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_908_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp532x_xop_905,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_53_909,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_928_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_928_inst_req_0;
      type_cast_928_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_928_inst_req_1;
      type_cast_928_inst_ack_1<= rack(0);
      type_cast_928_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_928_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext526_950,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_928_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_94_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_94_inst_req_0;
      type_cast_94_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_94_inst_req_1;
      type_cast_94_inst_ack_1<= rack(0);
      type_cast_94_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_94_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_91,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_95,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_972_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_972_inst_req_0;
      type_cast_972_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_972_inst_req_1;
      type_cast_972_inst_ack_1<= rack(0);
      type_cast_972_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_972_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_971_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv276_973,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1367_index_1_rename
    process(R_indvar_1366_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1366_resized;
      ov(13 downto 0) := iv;
      R_indvar_1366_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1367_index_1_resize
    process(indvar_1355) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1355;
      ov := iv(13 downto 0);
      R_indvar_1366_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1367_root_address_inst
    process(array_obj_ref_1367_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1367_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1367_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_486_index_1_rename
    process(R_indvar555_485_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar555_485_resized;
      ov(13 downto 0) := iv;
      R_indvar555_485_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_486_index_1_resize
    process(indvar555_474) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar555_474;
      ov := iv(13 downto 0);
      R_indvar555_485_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_486_root_address_inst
    process(array_obj_ref_486_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_486_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_486_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_693_index_1_rename
    process(R_indvar539_692_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar539_692_resized;
      ov(10 downto 0) := iv;
      R_indvar539_692_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_693_index_1_resize
    process(indvar539_681) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar539_681;
      ov := iv(10 downto 0);
      R_indvar539_692_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_693_root_address_inst
    process(array_obj_ref_693_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_693_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_693_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_937_index_1_rename
    process(R_indvar525_936_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar525_936_resized;
      ov(13 downto 0) := iv;
      R_indvar525_936_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_937_index_1_resize
    process(indvar525_925) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar525_925;
      ov := iv(13 downto 0);
      R_indvar525_936_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_937_root_address_inst
    process(array_obj_ref_937_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_937_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_937_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1372_addr_0
    process(ptr_deref_1372_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1372_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1372_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1372_base_resize
    process(arrayidx432_1369) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx432_1369;
      ov := iv(13 downto 0);
      ptr_deref_1372_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1372_gather_scatter
    process(ptr_deref_1372_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1372_data_0;
      ov(63 downto 0) := iv;
      tmp433_1373 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1372_root_address_inst
    process(ptr_deref_1372_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1372_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1372_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_623_addr_0
    process(ptr_deref_623_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_623_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_623_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_623_base_resize
    process(arrayidx_488) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_488;
      ov := iv(13 downto 0);
      ptr_deref_623_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_623_gather_scatter
    process(add186_621) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add186_621;
      ov(63 downto 0) := iv;
      ptr_deref_623_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_623_root_address_inst
    process(ptr_deref_623_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_623_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_623_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_830_addr_0
    process(ptr_deref_830_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_830_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_830_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_830_base_resize
    process(arrayidx246_695) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx246_695;
      ov := iv(10 downto 0);
      ptr_deref_830_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_830_gather_scatter
    process(add242_828) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add242_828;
      ov(63 downto 0) := iv;
      ptr_deref_830_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_830_root_address_inst
    process(ptr_deref_830_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_830_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_830_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_941_addr_0
    process(ptr_deref_941_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_941_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_941_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_941_base_resize
    process(arrayidx269_939) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx269_939;
      ov := iv(13 downto 0);
      ptr_deref_941_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_941_gather_scatter
    process(type_cast_943_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_943_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_941_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_941_root_address_inst
    process(ptr_deref_941_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_941_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_941_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1311_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264505_880;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1311_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1311_branch_req_0,
          ack0 => if_stmt_1311_branch_ack_0,
          ack1 => if_stmt_1311_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1483_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1482;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1483_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1483_branch_req_0,
          ack0 => if_stmt_1483_branch_ack_0,
          ack1 => if_stmt_1483_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_421_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp513_420;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_421_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_421_branch_req_0,
          ack0 => if_stmt_421_branch_ack_0,
          ack1 => if_stmt_421_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_436_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp194509_435;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_436_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_436_branch_req_0,
          ack0 => if_stmt_436_branch_ack_0,
          ack1 => if_stmt_436_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_637_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_636;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_637_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_637_branch_req_0,
          ack0 => if_stmt_637_branch_ack_0,
          ack1 => if_stmt_637_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_844_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_843;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_844_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_844_branch_req_0,
          ack0 => if_stmt_844_branch_ack_0,
          ack1 => if_stmt_844_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_881_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264505_880;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_881_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_881_branch_req_0,
          ack0 => if_stmt_881_branch_ack_0,
          ack1 => if_stmt_881_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_956_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_955;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_956_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_956_branch_req_0,
          ack0 => if_stmt_956_branch_ack_0,
          ack1 => if_stmt_956_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1334_inst
    process(tmp520_1323) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp520_1323, type_cast_1333_wire_constant, tmp_var);
      tmp520x_xop_1335 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_257_inst
    process(add74_253, shr_241) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add74_253, shr_241, tmp_var);
      add79_258 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_453_inst
    process(shr_241) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr_241, type_cast_452_wire_constant, tmp_var);
      tmp562x_xop_454 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_660_inst
    process(tmp548_649) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp548_649, type_cast_659_wire_constant, tmp_var);
      tmp548x_xop_661 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_904_inst
    process(tmp532_893) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp532_893, type_cast_903_wire_constant, tmp_var);
      tmp532x_xop_905 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1344_inst
    process(iNsTr_195_1339) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_195_1339, type_cast_1343_wire_constant, tmp_var);
      xx_xop_1345 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1476_inst
    process(indvar_1355) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1355, type_cast_1475_wire_constant, tmp_var);
      indvarx_xnext_1477 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_463_inst
    process(iNsTr_26_458) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_26_458, type_cast_462_wire_constant, tmp_var);
      xx_xop571_464 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_630_inst
    process(indvar555_474) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar555_474, type_cast_629_wire_constant, tmp_var);
      indvarx_xnext556_631 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_670_inst
    process(iNsTr_39_665) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_39_665, type_cast_669_wire_constant, tmp_var);
      xx_xop570_671 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_837_inst
    process(indvar539_681) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar539_681, type_cast_836_wire_constant, tmp_var);
      indvarx_xnext540_838 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_914_inst
    process(iNsTr_53_909) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_53_909, type_cast_913_wire_constant, tmp_var);
      xx_xop569_915 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_949_inst
    process(indvar525_925) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar525_925, type_cast_948_wire_constant, tmp_var);
      indvarx_xnext526_950 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_252_inst
    process(iNsTr_14_247) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_14_247, type_cast_251_wire_constant, tmp_var);
      add74_253 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1481_inst
    process(indvarx_xnext_1477, tmp524_1352) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1477, tmp524_1352, tmp_var);
      exitcond1_1482 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_635_inst
    process(indvarx_xnext556_631, tmp567_471) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext556_631, tmp567_471, tmp_var);
      exitcond3_636 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_842_inst
    process(indvarx_xnext540_838, tmp553_678) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext540_838, tmp553_678, tmp_var);
      exitcond2_843 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_954_inst
    process(indvarx_xnext526_950, tmp537_922) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext526_950, tmp537_922, tmp_var);
      exitcond_955 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1050_inst
    process(mul66_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_235, type_cast_1049_wire_constant, tmp_var);
      shr304_1051 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1106_inst
    process(mul66_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_235, type_cast_1105_wire_constant, tmp_var);
      shr321_1107 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1162_inst
    process(add79_258) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_258, type_cast_1161_wire_constant, tmp_var);
      shr338_1163 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1322_inst
    process(mul259_874) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_874, type_cast_1321_wire_constant, tmp_var);
      tmp520_1323 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_240_inst
    process(mul66_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_235, type_cast_239_wire_constant, tmp_var);
      shr_241 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_246_inst
    process(mul66_235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_235, type_cast_245_wire_constant, tmp_var);
      iNsTr_14_247 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_648_inst
    process(mul91_289) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul91_289, type_cast_647_wire_constant, tmp_var);
      tmp548_649 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_892_inst
    process(mul259_874) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_874, type_cast_891_wire_constant, tmp_var);
      tmp532_893 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1220_inst
    process(sub_1211) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1211, type_cast_1219_wire_constant, tmp_var);
      shr364_1221 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1230_inst
    process(sub_1211) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1211, type_cast_1229_wire_constant, tmp_var);
      shr370_1231 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1240_inst
    process(sub_1211) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1211, type_cast_1239_wire_constant, tmp_var);
      shr376_1241 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1250_inst
    process(sub_1211) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1211, type_cast_1249_wire_constant, tmp_var);
      shr382_1251 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1260_inst
    process(sub_1211) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1211, type_cast_1259_wire_constant, tmp_var);
      shr388_1261 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1270_inst
    process(sub_1211) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1211, type_cast_1269_wire_constant, tmp_var);
      shr394_1271 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1280_inst
    process(sub_1211) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1211, type_cast_1279_wire_constant, tmp_var);
      shr400_1281 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1382_inst
    process(tmp433_1373) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1373, type_cast_1381_wire_constant, tmp_var);
      shr440_1383 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1392_inst
    process(tmp433_1373) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1373, type_cast_1391_wire_constant, tmp_var);
      shr446_1393 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1402_inst
    process(tmp433_1373) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1373, type_cast_1401_wire_constant, tmp_var);
      shr452_1403 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1412_inst
    process(tmp433_1373) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1373, type_cast_1411_wire_constant, tmp_var);
      shr458_1413 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1422_inst
    process(tmp433_1373) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1373, type_cast_1421_wire_constant, tmp_var);
      shr464_1423 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1432_inst
    process(tmp433_1373) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1373, type_cast_1431_wire_constant, tmp_var);
      shr470_1433 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1442_inst
    process(tmp433_1373) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp433_1373, type_cast_1441_wire_constant, tmp_var);
      shr476_1443 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_229_inst
    process(conv63_221, conv61_217) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv63_221, conv61_217, tmp_var);
      mul_230 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_234_inst
    process(mul_230, conv65_225) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_230, conv65_225, tmp_var);
      mul66_235 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_278_inst
    process(conv84_266, conv82_262) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv84_266, conv82_262, tmp_var);
      mul85_279 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_283_inst
    process(mul85_279, conv87_270) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul85_279, conv87_270, tmp_var);
      mul88_284 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_288_inst
    process(mul88_284, conv90_274) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul88_284, conv90_274, tmp_var);
      mul91_289 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_868_inst
    process(conv255_860, conv253_856) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv255_860, conv253_856, tmp_var);
      mul256_869 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_873_inst
    process(mul256_869, conv258_864) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul256_869, conv258_864, tmp_var);
      mul259_874 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_112_inst
    process(shl18_101, conv20_108) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_101, conv20_108, tmp_var);
      add21_113 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_137_inst
    process(shl27_126, conv29_133) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_126, conv29_133, tmp_var);
      add30_138 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_162_inst
    process(shl36_151, conv38_158) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_151, conv38_158, tmp_var);
      add39_163 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_187_inst
    process(shl45_176, conv47_183) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_176, conv47_183, tmp_var);
      add48_188 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_212_inst
    process(shl54_201, conv56_208) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_201, conv56_208, tmp_var);
      add57_213 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_313_inst
    process(shl96_302, conv98_309) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl96_302, conv98_309, tmp_var);
      add99_314 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_338_inst
    process(shl105_327, conv107_334) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_327, conv107_334, tmp_var);
      add108_339 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_363_inst
    process(shl114_352, conv116_359) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_352, conv116_359, tmp_var);
      add117_364 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_388_inst
    process(shl123_377, conv125_384) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl123_377, conv125_384, tmp_var);
      add126_389 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_413_inst
    process(shl132_402, conv134_409) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_402, conv134_409, tmp_var);
      add135_414 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_62_inst
    process(shl_51, conv3_58) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_51, conv3_58, tmp_var);
      add_63 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_87_inst
    process(shl9_76, conv11_83) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_76, conv11_83, tmp_var);
      add12_88 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_512_inst
    process(shl146_501, conv149_508) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl146_501, conv149_508, tmp_var);
      add150_513 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_530_inst
    process(shl152_519, conv155_526) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl152_519, conv155_526, tmp_var);
      add156_531 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_548_inst
    process(shl158_537, conv161_544) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl158_537, conv161_544, tmp_var);
      add162_549 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_566_inst
    process(shl164_555, conv167_562) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl164_555, conv167_562, tmp_var);
      add168_567 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_584_inst
    process(shl170_573, conv173_580) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl170_573, conv173_580, tmp_var);
      add174_585 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_602_inst
    process(shl176_591, conv179_598) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl176_591, conv179_598, tmp_var);
      add180_603 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_620_inst
    process(shl182_609, conv185_616) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl182_609, conv185_616, tmp_var);
      add186_621 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_719_inst
    process(shl202_708, conv205_715) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl202_708, conv205_715, tmp_var);
      add206_720 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_737_inst
    process(shl208_726, conv211_733) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl208_726, conv211_733, tmp_var);
      add212_738 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_755_inst
    process(shl214_744, conv217_751) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl214_744, conv217_751, tmp_var);
      add218_756 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_773_inst
    process(shl220_762, conv223_769) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl220_762, conv223_769, tmp_var);
      add224_774 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_791_inst
    process(shl226_780, conv229_787) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl226_780, conv229_787, tmp_var);
      add230_792 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_809_inst
    process(shl232_798, conv235_805) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl232_798, conv235_805, tmp_var);
      add236_810 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_827_inst
    process(shl238_816, conv241_823) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl238_816, conv241_823, tmp_var);
      add242_828 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_100_inst
    process(conv17_95) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_95, type_cast_99_wire_constant, tmp_var);
      shl18_101 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_125_inst
    process(conv26_120) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_120, type_cast_124_wire_constant, tmp_var);
      shl27_126 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_150_inst
    process(conv35_145) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_145, type_cast_149_wire_constant, tmp_var);
      shl36_151 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_175_inst
    process(conv44_170) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_170, type_cast_174_wire_constant, tmp_var);
      shl45_176 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_200_inst
    process(conv53_195) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_195, type_cast_199_wire_constant, tmp_var);
      shl54_201 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_301_inst
    process(conv95_296) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv95_296, type_cast_300_wire_constant, tmp_var);
      shl96_302 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_326_inst
    process(conv104_321) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv104_321, type_cast_325_wire_constant, tmp_var);
      shl105_327 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_351_inst
    process(conv113_346) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv113_346, type_cast_350_wire_constant, tmp_var);
      shl114_352 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_376_inst
    process(conv122_371) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv122_371, type_cast_375_wire_constant, tmp_var);
      shl123_377 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_401_inst
    process(conv131_396) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_396, type_cast_400_wire_constant, tmp_var);
      shl132_402 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_50_inst
    process(conv1_45) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_45, type_cast_49_wire_constant, tmp_var);
      shl_51 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_75_inst
    process(conv8_70) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_70, type_cast_74_wire_constant, tmp_var);
      shl9_76 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_500_inst
    process(conv144_495) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv144_495, type_cast_499_wire_constant, tmp_var);
      shl146_501 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_518_inst
    process(add150_513) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add150_513, type_cast_517_wire_constant, tmp_var);
      shl152_519 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_536_inst
    process(add156_531) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add156_531, type_cast_535_wire_constant, tmp_var);
      shl158_537 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_554_inst
    process(add162_549) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add162_549, type_cast_553_wire_constant, tmp_var);
      shl164_555 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_572_inst
    process(add168_567) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add168_567, type_cast_571_wire_constant, tmp_var);
      shl170_573 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_590_inst
    process(add174_585) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add174_585, type_cast_589_wire_constant, tmp_var);
      shl176_591 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_608_inst
    process(add180_603) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add180_603, type_cast_607_wire_constant, tmp_var);
      shl182_609 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_707_inst
    process(conv200_702) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv200_702, type_cast_706_wire_constant, tmp_var);
      shl202_708 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_725_inst
    process(add206_720) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add206_720, type_cast_724_wire_constant, tmp_var);
      shl208_726 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_743_inst
    process(add212_738) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add212_738, type_cast_742_wire_constant, tmp_var);
      shl214_744 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_761_inst
    process(add218_756) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add218_756, type_cast_760_wire_constant, tmp_var);
      shl220_762 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_779_inst
    process(add224_774) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add224_774, type_cast_778_wire_constant, tmp_var);
      shl226_780 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_797_inst
    process(add230_792) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add230_792, type_cast_796_wire_constant, tmp_var);
      shl232_798 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_815_inst
    process(add236_810) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add236_810, type_cast_814_wire_constant, tmp_var);
      shl238_816 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1210_inst
    process(conv355_1206, conv276_973) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv355_1206, conv276_973, tmp_var);
      sub_1211 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1328_inst
    process(tmp520_1323) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp520_1323, type_cast_1327_wire_constant, tmp_var);
      tmp521_1329 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_419_inst
    process(mul66_235) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul66_235, type_cast_418_wire_constant, tmp_var);
      cmp513_420 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_434_inst
    process(mul91_289) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul91_289, type_cast_433_wire_constant, tmp_var);
      cmp194509_435 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_447_inst
    process(shr_241) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_241, type_cast_446_wire_constant, tmp_var);
      tmp563_448 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_654_inst
    process(tmp548_649) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp548_649, type_cast_653_wire_constant, tmp_var);
      tmp549_655 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_879_inst
    process(mul259_874) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul259_874, type_cast_878_wire_constant, tmp_var);
      cmp264505_880 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_898_inst
    process(tmp532_893) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp532_893, type_cast_897_wire_constant, tmp_var);
      tmp533_899 <= tmp_var; --
    end process;
    -- shared split operator group (107) : array_obj_ref_1367_index_offset 
    ApIntAdd_group_107: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1366_scaled;
      array_obj_ref_1367_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1367_index_offset_req_0;
      array_obj_ref_1367_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1367_index_offset_req_1;
      array_obj_ref_1367_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_107_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_107_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_107",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 107
    -- shared split operator group (108) : array_obj_ref_486_index_offset 
    ApIntAdd_group_108: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar555_485_scaled;
      array_obj_ref_486_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_486_index_offset_req_0;
      array_obj_ref_486_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_486_index_offset_req_1;
      array_obj_ref_486_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_108_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_108_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_108",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 108
    -- shared split operator group (109) : array_obj_ref_693_index_offset 
    ApIntAdd_group_109: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar539_692_scaled;
      array_obj_ref_693_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_693_index_offset_req_0;
      array_obj_ref_693_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_693_index_offset_req_1;
      array_obj_ref_693_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_109_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_109_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_109",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100010",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 109
    -- shared split operator group (110) : array_obj_ref_937_index_offset 
    ApIntAdd_group_110: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar525_936_scaled;
      array_obj_ref_937_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_937_index_offset_req_0;
      array_obj_ref_937_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_937_index_offset_req_1;
      array_obj_ref_937_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_110_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_110_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_110",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 110
    -- unary operator type_cast_1204_inst
    process(call354_1201) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call354_1201, tmp_var);
      type_cast_1204_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_971_inst
    process(call275_967) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call275_967, tmp_var);
      type_cast_971_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1372_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1372_load_0_req_0;
      ptr_deref_1372_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1372_load_0_req_1;
      ptr_deref_1372_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1372_word_address_0;
      ptr_deref_1372_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(13 downto 0),
          mtag => memory_space_2_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_623_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_623_store_0_req_0;
      ptr_deref_623_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_623_store_0_req_1;
      ptr_deref_623_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_623_word_address_0;
      data_in <= ptr_deref_623_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_830_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_830_store_0_req_0;
      ptr_deref_830_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_830_store_0_req_1;
      ptr_deref_830_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_830_word_address_0;
      data_in <= ptr_deref_830_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(10 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_941_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_941_store_0_req_0;
      ptr_deref_941_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_941_store_0_req_1;
      ptr_deref_941_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_941_word_address_0;
      data_in <= ptr_deref_941_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Block0_done_1188_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1188_inst_req_0;
      RPIPE_Block0_done_1188_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1188_inst_req_1;
      RPIPE_Block0_done_1188_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call346_1189 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1191_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1191_inst_req_0;
      RPIPE_Block1_done_1191_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1191_inst_req_1;
      RPIPE_Block1_done_1191_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call348_1192 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1194_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1194_inst_req_0;
      RPIPE_Block2_done_1194_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1194_inst_req_1;
      RPIPE_Block2_done_1194_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call350_1195 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1197_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1197_inst_req_0;
      RPIPE_Block3_done_1197_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1197_inst_req_1;
      RPIPE_Block3_done_1197_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call352_1198 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_ConvTranspose_input_pipe_710_inst RPIPE_ConvTranspose_input_pipe_53_inst RPIPE_ConvTranspose_input_pipe_128_inst RPIPE_ConvTranspose_input_pipe_40_inst RPIPE_ConvTranspose_input_pipe_782_inst RPIPE_ConvTranspose_input_pipe_153_inst RPIPE_ConvTranspose_input_pipe_800_inst RPIPE_ConvTranspose_input_pipe_165_inst RPIPE_ConvTranspose_input_pipe_140_inst RPIPE_ConvTranspose_input_pipe_190_inst RPIPE_ConvTranspose_input_pipe_78_inst RPIPE_ConvTranspose_input_pipe_115_inst RPIPE_ConvTranspose_input_pipe_728_inst RPIPE_ConvTranspose_input_pipe_178_inst RPIPE_ConvTranspose_input_pipe_818_inst RPIPE_ConvTranspose_input_pipe_746_inst RPIPE_ConvTranspose_input_pipe_697_inst RPIPE_ConvTranspose_input_pipe_764_inst RPIPE_ConvTranspose_input_pipe_90_inst RPIPE_ConvTranspose_input_pipe_103_inst RPIPE_ConvTranspose_input_pipe_65_inst RPIPE_ConvTranspose_input_pipe_203_inst RPIPE_ConvTranspose_input_pipe_291_inst RPIPE_ConvTranspose_input_pipe_304_inst RPIPE_ConvTranspose_input_pipe_316_inst RPIPE_ConvTranspose_input_pipe_329_inst RPIPE_ConvTranspose_input_pipe_341_inst RPIPE_ConvTranspose_input_pipe_354_inst RPIPE_ConvTranspose_input_pipe_366_inst RPIPE_ConvTranspose_input_pipe_379_inst RPIPE_ConvTranspose_input_pipe_391_inst RPIPE_ConvTranspose_input_pipe_404_inst RPIPE_ConvTranspose_input_pipe_490_inst RPIPE_ConvTranspose_input_pipe_503_inst RPIPE_ConvTranspose_input_pipe_521_inst RPIPE_ConvTranspose_input_pipe_539_inst RPIPE_ConvTranspose_input_pipe_557_inst RPIPE_ConvTranspose_input_pipe_575_inst RPIPE_ConvTranspose_input_pipe_593_inst RPIPE_ConvTranspose_input_pipe_611_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_710_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_53_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_128_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_40_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_782_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_153_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_800_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_165_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_140_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_190_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_78_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_115_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_728_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_178_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_818_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_746_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_697_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_764_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_90_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_103_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_65_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_203_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_291_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_304_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_316_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_329_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_341_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_354_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_366_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_379_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_391_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_404_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_490_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_503_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_521_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_539_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_557_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_575_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_593_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_611_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_710_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_53_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_128_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_40_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_782_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_153_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_800_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_165_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_140_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_190_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_78_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_115_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_728_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_178_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_818_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_746_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_697_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_764_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_90_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_103_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_65_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_203_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_291_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_304_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_316_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_329_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_341_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_354_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_366_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_379_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_391_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_404_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_490_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_503_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_521_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_539_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_557_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_575_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_593_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_611_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_710_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_53_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_128_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_40_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_782_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_153_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_800_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_165_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_140_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_190_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_78_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_115_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_728_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_178_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_818_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_746_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_697_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_764_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_90_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_103_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_65_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_203_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_291_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_304_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_316_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_329_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_341_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_354_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_366_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_379_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_391_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_404_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_490_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_503_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_521_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_539_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_557_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_575_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_593_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_611_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_710_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_53_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_128_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_40_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_782_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_153_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_800_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_165_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_140_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_190_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_78_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_115_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_728_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_178_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_818_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_746_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_697_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_764_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_90_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_103_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_65_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_203_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_291_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_304_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_316_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_329_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_341_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_354_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_366_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_379_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_391_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_404_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_490_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_503_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_521_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_539_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_557_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_575_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_593_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_611_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call203_711 <= data_out(319 downto 312);
      call2_54 <= data_out(311 downto 304);
      call28_129 <= data_out(303 downto 296);
      call_41 <= data_out(295 downto 288);
      call227_783 <= data_out(287 downto 280);
      call37_154 <= data_out(279 downto 272);
      call233_801 <= data_out(271 downto 264);
      call41_166 <= data_out(263 downto 256);
      call32_141 <= data_out(255 downto 248);
      call50_191 <= data_out(247 downto 240);
      call10_79 <= data_out(239 downto 232);
      call23_116 <= data_out(231 downto 224);
      call209_729 <= data_out(223 downto 216);
      call46_179 <= data_out(215 downto 208);
      call239_819 <= data_out(207 downto 200);
      call215_747 <= data_out(199 downto 192);
      call199_698 <= data_out(191 downto 184);
      call221_765 <= data_out(183 downto 176);
      call14_91 <= data_out(175 downto 168);
      call19_104 <= data_out(167 downto 160);
      call5_66 <= data_out(159 downto 152);
      call55_204 <= data_out(151 downto 144);
      call92_292 <= data_out(143 downto 136);
      call97_305 <= data_out(135 downto 128);
      call101_317 <= data_out(127 downto 120);
      call106_330 <= data_out(119 downto 112);
      call110_342 <= data_out(111 downto 104);
      call115_355 <= data_out(103 downto 96);
      call119_367 <= data_out(95 downto 88);
      call124_380 <= data_out(87 downto 80);
      call128_392 <= data_out(79 downto 72);
      call133_405 <= data_out(71 downto 64);
      call143_491 <= data_out(63 downto 56);
      call147_504 <= data_out(55 downto 48);
      call153_522 <= data_out(47 downto 40);
      call159_540 <= data_out(39 downto 32);
      call165_558 <= data_out(31 downto 24);
      call171_576 <= data_out(23 downto 16);
      call177_594 <= data_out(15 downto 8);
      call183_612 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_4_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_4: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_4", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_Block0_start_978_inst WPIPE_Block0_start_975_inst WPIPE_Block0_start_1010_inst WPIPE_Block0_start_1013_inst WPIPE_Block0_start_1016_inst WPIPE_Block0_start_999_inst WPIPE_Block0_start_981_inst WPIPE_Block0_start_984_inst WPIPE_Block0_start_987_inst WPIPE_Block0_start_1006_inst WPIPE_Block0_start_990_inst WPIPE_Block0_start_1002_inst WPIPE_Block0_start_993_inst WPIPE_Block0_start_996_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block0_start_978_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block0_start_975_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block0_start_1010_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block0_start_1013_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block0_start_1016_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block0_start_999_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block0_start_981_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block0_start_984_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_start_987_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_start_1006_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_start_990_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_start_1002_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_start_993_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_start_996_inst_req_0;
      WPIPE_Block0_start_978_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block0_start_975_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block0_start_1010_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block0_start_1013_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block0_start_1016_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block0_start_999_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block0_start_981_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block0_start_984_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_start_987_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_start_1006_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_start_990_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_start_1002_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_start_993_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_start_996_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block0_start_978_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block0_start_975_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block0_start_1010_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block0_start_1013_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block0_start_1016_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block0_start_999_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block0_start_981_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block0_start_984_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_start_987_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_start_1006_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_start_990_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_start_1002_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_start_993_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_start_996_inst_req_1;
      WPIPE_Block0_start_978_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block0_start_975_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block0_start_1010_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block0_start_1013_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block0_start_1016_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block0_start_999_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block0_start_981_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block0_start_984_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_start_987_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_start_1006_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_start_990_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_start_1002_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_start_993_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_start_996_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add12_88 & add_63 & add117_364 & add126_389 & add135_414 & add108_339 & add21_113 & add30_138 & add39_163 & type_cast_1008_wire_constant & add48_188 & type_cast_1004_wire_constant & add57_213 & add99_314;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1056_inst WPIPE_Block1_start_1072_inst WPIPE_Block1_start_1069_inst WPIPE_Block1_start_1066_inst WPIPE_Block1_start_1043_inst WPIPE_Block1_start_1019_inst WPIPE_Block1_start_1040_inst WPIPE_Block1_start_1022_inst WPIPE_Block1_start_1025_inst WPIPE_Block1_start_1063_inst WPIPE_Block1_start_1028_inst WPIPE_Block1_start_1031_inst WPIPE_Block1_start_1034_inst WPIPE_Block1_start_1037_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block1_start_1056_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block1_start_1072_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block1_start_1069_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block1_start_1066_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block1_start_1043_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block1_start_1019_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block1_start_1040_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block1_start_1022_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block1_start_1025_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block1_start_1063_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block1_start_1028_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block1_start_1031_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block1_start_1034_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block1_start_1037_inst_req_0;
      WPIPE_Block1_start_1056_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block1_start_1072_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block1_start_1069_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block1_start_1066_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block1_start_1043_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block1_start_1019_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block1_start_1040_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block1_start_1022_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block1_start_1025_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block1_start_1063_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block1_start_1028_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block1_start_1031_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block1_start_1034_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block1_start_1037_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block1_start_1056_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block1_start_1072_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block1_start_1069_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block1_start_1066_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block1_start_1043_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block1_start_1019_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block1_start_1040_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block1_start_1022_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block1_start_1025_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block1_start_1063_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block1_start_1028_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block1_start_1031_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block1_start_1034_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block1_start_1037_inst_req_1;
      WPIPE_Block1_start_1056_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block1_start_1072_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block1_start_1069_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block1_start_1066_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block1_start_1043_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block1_start_1019_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block1_start_1040_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block1_start_1022_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block1_start_1025_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block1_start_1063_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block1_start_1028_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block1_start_1031_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block1_start_1034_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block1_start_1037_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= conv305_1055 & add135_414 & add126_389 & add117_364 & add108_339 & add_63 & add99_314 & add12_88 & add21_113 & conv307_1062 & add30_138 & add39_163 & add48_188 & add57_213;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1125_inst WPIPE_Block2_start_1081_inst WPIPE_Block2_start_1078_inst WPIPE_Block2_start_1075_inst WPIPE_Block2_start_1084_inst WPIPE_Block2_start_1128_inst WPIPE_Block2_start_1087_inst WPIPE_Block2_start_1090_inst WPIPE_Block2_start_1093_inst WPIPE_Block2_start_1096_inst WPIPE_Block2_start_1099_inst WPIPE_Block2_start_1112_inst WPIPE_Block2_start_1119_inst WPIPE_Block2_start_1122_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block2_start_1125_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block2_start_1081_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block2_start_1078_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block2_start_1075_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block2_start_1084_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block2_start_1128_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block2_start_1087_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block2_start_1090_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block2_start_1093_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block2_start_1096_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block2_start_1099_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block2_start_1112_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block2_start_1119_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block2_start_1122_inst_req_0;
      WPIPE_Block2_start_1125_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block2_start_1081_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block2_start_1078_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block2_start_1075_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block2_start_1084_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block2_start_1128_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block2_start_1087_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block2_start_1090_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block2_start_1093_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block2_start_1096_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block2_start_1099_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block2_start_1112_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block2_start_1119_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block2_start_1122_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block2_start_1125_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block2_start_1081_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block2_start_1078_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block2_start_1075_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block2_start_1084_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block2_start_1128_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block2_start_1087_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block2_start_1090_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block2_start_1093_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block2_start_1096_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block2_start_1099_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block2_start_1112_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block2_start_1119_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block2_start_1122_inst_req_1;
      WPIPE_Block2_start_1125_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block2_start_1081_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block2_start_1078_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block2_start_1075_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block2_start_1084_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block2_start_1128_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block2_start_1087_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block2_start_1090_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block2_start_1093_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block2_start_1096_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block2_start_1099_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block2_start_1112_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block2_start_1119_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block2_start_1122_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add126_389 & add21_113 & add12_88 & add_63 & add30_138 & add135_414 & add39_163 & add48_188 & add57_213 & add99_314 & add108_339 & conv322_1111 & conv324_1118 & add117_364;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1155_inst WPIPE_Block3_start_1181_inst WPIPE_Block3_start_1131_inst WPIPE_Block3_start_1134_inst WPIPE_Block3_start_1146_inst WPIPE_Block3_start_1184_inst WPIPE_Block3_start_1152_inst WPIPE_Block3_start_1149_inst WPIPE_Block3_start_1175_inst WPIPE_Block3_start_1168_inst WPIPE_Block3_start_1178_inst WPIPE_Block3_start_1140_inst WPIPE_Block3_start_1137_inst WPIPE_Block3_start_1143_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(223 downto 0);
      signal sample_req, sample_ack : BooleanArray( 13 downto 0);
      signal update_req, update_ack : BooleanArray( 13 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 13 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant inBUFs : IntegerArray(13 downto 0) := (13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      sample_req_unguarded(13) <= WPIPE_Block3_start_1155_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Block3_start_1181_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block3_start_1131_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block3_start_1134_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block3_start_1146_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block3_start_1184_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block3_start_1152_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block3_start_1149_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block3_start_1175_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block3_start_1168_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block3_start_1178_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block3_start_1140_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block3_start_1137_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block3_start_1143_inst_req_0;
      WPIPE_Block3_start_1155_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Block3_start_1181_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block3_start_1131_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block3_start_1134_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block3_start_1146_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block3_start_1184_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block3_start_1152_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block3_start_1149_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block3_start_1175_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block3_start_1168_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block3_start_1178_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block3_start_1140_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block3_start_1137_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block3_start_1143_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(13) <= WPIPE_Block3_start_1155_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Block3_start_1181_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block3_start_1131_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block3_start_1134_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block3_start_1146_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block3_start_1184_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block3_start_1152_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block3_start_1149_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block3_start_1175_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block3_start_1168_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block3_start_1178_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block3_start_1140_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block3_start_1137_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block3_start_1143_inst_req_1;
      WPIPE_Block3_start_1155_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Block3_start_1181_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block3_start_1131_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block3_start_1134_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block3_start_1146_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block3_start_1184_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block3_start_1152_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block3_start_1149_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block3_start_1175_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block3_start_1168_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block3_start_1178_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block3_start_1140_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block3_start_1137_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block3_start_1143_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      data_in <= add108_339 & add126_389 & add_63 & add12_88 & add48_188 & add135_414 & add99_314 & add57_213 & conv341_1174 & conv339_1167 & add117_364 & add30_138 & add21_113 & add39_163;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 14, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_ConvTranspose_output_pipe_1295_inst WPIPE_ConvTranspose_output_pipe_1307_inst WPIPE_ConvTranspose_output_pipe_1301_inst WPIPE_ConvTranspose_output_pipe_1298_inst WPIPE_ConvTranspose_output_pipe_1304_inst WPIPE_ConvTranspose_output_pipe_1286_inst WPIPE_ConvTranspose_output_pipe_1289_inst WPIPE_ConvTranspose_output_pipe_1292_inst WPIPE_ConvTranspose_output_pipe_1448_inst WPIPE_ConvTranspose_output_pipe_1451_inst WPIPE_ConvTranspose_output_pipe_1454_inst WPIPE_ConvTranspose_output_pipe_1457_inst WPIPE_ConvTranspose_output_pipe_1460_inst WPIPE_ConvTranspose_output_pipe_1463_inst WPIPE_ConvTranspose_output_pipe_1466_inst WPIPE_ConvTranspose_output_pipe_1469_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 15 downto 0);
      signal update_req, update_ack : BooleanArray( 15 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 15 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      sample_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1295_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1307_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1301_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1298_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1304_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1286_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1289_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1292_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1448_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1451_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1454_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1457_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1460_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1463_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1466_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1469_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1295_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1307_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1301_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1298_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1304_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1286_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1289_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1292_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1448_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1451_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1454_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1457_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1460_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1463_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1466_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1469_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(15) <= WPIPE_ConvTranspose_output_pipe_1295_inst_req_1;
      update_req_unguarded(14) <= WPIPE_ConvTranspose_output_pipe_1307_inst_req_1;
      update_req_unguarded(13) <= WPIPE_ConvTranspose_output_pipe_1301_inst_req_1;
      update_req_unguarded(12) <= WPIPE_ConvTranspose_output_pipe_1298_inst_req_1;
      update_req_unguarded(11) <= WPIPE_ConvTranspose_output_pipe_1304_inst_req_1;
      update_req_unguarded(10) <= WPIPE_ConvTranspose_output_pipe_1286_inst_req_1;
      update_req_unguarded(9) <= WPIPE_ConvTranspose_output_pipe_1289_inst_req_1;
      update_req_unguarded(8) <= WPIPE_ConvTranspose_output_pipe_1292_inst_req_1;
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1448_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1451_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1454_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1457_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1460_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1463_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1466_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1469_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1295_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_ConvTranspose_output_pipe_1307_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_ConvTranspose_output_pipe_1301_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_ConvTranspose_output_pipe_1298_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_ConvTranspose_output_pipe_1304_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_ConvTranspose_output_pipe_1286_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_ConvTranspose_output_pipe_1289_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_ConvTranspose_output_pipe_1292_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_ConvTranspose_output_pipe_1448_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1451_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1454_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1457_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1460_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1463_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1466_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1469_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      data_in <= conv385_1255 & conv361_1215 & conv373_1235 & conv379_1245 & conv367_1225 & conv403_1285 & conv397_1275 & conv391_1265 & conv479_1447 & conv473_1437 & conv467_1427 & conv461_1417 & conv455_1407 & conv449_1397 & conv443_1387 & conv437_1377;
      ConvTranspose_output_pipe_write_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_4_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 16, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared call operator group (0) : call_stmt_967_call call_stmt_1201_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_967_call_req_0;
      reqL_unguarded(0) <= call_stmt_1201_call_req_0;
      call_stmt_967_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1201_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_967_call_req_1;
      reqR_unguarded(0) <= call_stmt_1201_call_req_1;
      call_stmt_967_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1201_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call275_967 <= data_out(127 downto 64);
      call354_1201 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3758_start: Boolean;
  signal convTransposeA_CP_3758_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block0_start_1514_inst_req_1 : boolean;
  signal phi_stmt_1627_ack_0 : boolean;
  signal RPIPE_Block0_start_1517_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1517_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1499_inst_ack_0 : boolean;
  signal phi_stmt_1606_ack_0 : boolean;
  signal RPIPE_Block0_start_1511_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1520_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1499_inst_req_0 : boolean;
  signal type_cast_1543_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1511_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1508_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1505_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1505_inst_ack_1 : boolean;
  signal type_cast_1633_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1557_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1557_inst_ack_1 : boolean;
  signal phi_stmt_1620_ack_0 : boolean;
  signal RPIPE_Block0_start_1502_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1520_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1505_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1502_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1505_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1514_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1554_inst_req_0 : boolean;
  signal phi_stmt_1822_ack_0 : boolean;
  signal type_cast_1543_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1554_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1517_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1517_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1523_inst_ack_0 : boolean;
  signal type_cast_1530_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1557_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1523_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1523_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1514_inst_ack_1 : boolean;
  signal phi_stmt_1627_req_1 : boolean;
  signal RPIPE_Block0_start_1514_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1511_inst_ack_0 : boolean;
  signal type_cast_1530_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1508_inst_ack_0 : boolean;
  signal type_cast_1612_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1511_inst_req_1 : boolean;
  signal phi_stmt_1613_ack_0 : boolean;
  signal RPIPE_Block0_start_1523_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1557_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1539_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1508_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1502_inst_req_0 : boolean;
  signal type_cast_1530_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1508_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1554_inst_ack_0 : boolean;
  signal type_cast_1543_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1539_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1499_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1499_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1539_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1539_inst_ack_0 : boolean;
  signal type_cast_1530_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1502_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1554_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1520_inst_req_0 : boolean;
  signal type_cast_1633_inst_ack_1 : boolean;
  signal type_cast_1543_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1520_inst_ack_0 : boolean;
  signal phi_stmt_1606_req_0 : boolean;
  signal type_cast_1588_inst_req_1 : boolean;
  signal phi_stmt_1815_req_0 : boolean;
  signal type_cast_1588_inst_ack_1 : boolean;
  signal type_cast_1592_inst_req_0 : boolean;
  signal type_cast_1592_inst_ack_0 : boolean;
  signal type_cast_1588_inst_ack_0 : boolean;
  signal type_cast_1588_inst_req_0 : boolean;
  signal type_cast_1633_inst_req_0 : boolean;
  signal type_cast_1821_inst_ack_1 : boolean;
  signal type_cast_1821_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1551_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1526_inst_ack_1 : boolean;
  signal type_cast_1584_inst_req_1 : boolean;
  signal type_cast_1584_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1551_inst_req_1 : boolean;
  signal phi_stmt_1815_ack_0 : boolean;
  signal RPIPE_Block0_start_1526_inst_req_1 : boolean;
  signal type_cast_1584_inst_ack_0 : boolean;
  signal phi_stmt_1815_req_1 : boolean;
  signal type_cast_1584_inst_req_0 : boolean;
  signal phi_stmt_1627_req_0 : boolean;
  signal type_cast_1633_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1551_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1526_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1551_inst_req_0 : boolean;
  signal type_cast_1592_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1526_inst_req_0 : boolean;
  signal type_cast_1592_inst_ack_1 : boolean;
  signal phi_stmt_1613_req_0 : boolean;
  signal type_cast_1821_inst_ack_0 : boolean;
  signal type_cast_1821_inst_req_0 : boolean;
  signal type_cast_1596_inst_req_0 : boolean;
  signal type_cast_1596_inst_ack_0 : boolean;
  signal type_cast_1596_inst_req_1 : boolean;
  signal type_cast_1596_inst_ack_1 : boolean;
  signal type_cast_1668_inst_req_0 : boolean;
  signal type_cast_1668_inst_ack_0 : boolean;
  signal type_cast_1668_inst_req_1 : boolean;
  signal type_cast_1668_inst_ack_1 : boolean;
  signal type_cast_1672_inst_req_0 : boolean;
  signal phi_stmt_1822_req_0 : boolean;
  signal type_cast_1672_inst_ack_0 : boolean;
  signal type_cast_1672_inst_req_1 : boolean;
  signal type_cast_1825_inst_ack_1 : boolean;
  signal type_cast_1672_inst_ack_1 : boolean;
  signal type_cast_1676_inst_req_0 : boolean;
  signal type_cast_1825_inst_req_1 : boolean;
  signal type_cast_1676_inst_ack_0 : boolean;
  signal type_cast_1676_inst_req_1 : boolean;
  signal type_cast_1676_inst_ack_1 : boolean;
  signal type_cast_1706_inst_req_0 : boolean;
  signal type_cast_1706_inst_ack_0 : boolean;
  signal type_cast_1706_inst_req_1 : boolean;
  signal type_cast_1825_inst_ack_0 : boolean;
  signal type_cast_1706_inst_ack_1 : boolean;
  signal phi_stmt_1822_req_1 : boolean;
  signal type_cast_1827_inst_ack_1 : boolean;
  signal type_cast_1827_inst_req_1 : boolean;
  signal type_cast_1827_inst_ack_0 : boolean;
  signal type_cast_1827_inst_req_0 : boolean;
  signal phi_stmt_1620_req_1 : boolean;
  signal type_cast_1626_inst_ack_1 : boolean;
  signal type_cast_1626_inst_req_1 : boolean;
  signal array_obj_ref_1712_index_offset_req_0 : boolean;
  signal type_cast_1825_inst_req_0 : boolean;
  signal array_obj_ref_1712_index_offset_ack_0 : boolean;
  signal array_obj_ref_1712_index_offset_req_1 : boolean;
  signal array_obj_ref_1712_index_offset_ack_1 : boolean;
  signal phi_stmt_1828_ack_0 : boolean;
  signal addr_of_1713_final_reg_req_0 : boolean;
  signal addr_of_1713_final_reg_ack_0 : boolean;
  signal addr_of_1713_final_reg_req_1 : boolean;
  signal addr_of_1713_final_reg_ack_1 : boolean;
  signal type_cast_1626_inst_ack_0 : boolean;
  signal type_cast_1626_inst_req_0 : boolean;
  signal phi_stmt_1606_req_1 : boolean;
  signal type_cast_1612_inst_ack_1 : boolean;
  signal ptr_deref_1717_load_0_req_0 : boolean;
  signal ptr_deref_1717_load_0_ack_0 : boolean;
  signal type_cast_1612_inst_req_1 : boolean;
  signal ptr_deref_1717_load_0_req_1 : boolean;
  signal ptr_deref_1717_load_0_ack_1 : boolean;
  signal phi_stmt_1828_req_0 : boolean;
  signal type_cast_1831_inst_ack_1 : boolean;
  signal type_cast_1831_inst_req_1 : boolean;
  signal array_obj_ref_1735_index_offset_req_0 : boolean;
  signal array_obj_ref_1735_index_offset_ack_0 : boolean;
  signal array_obj_ref_1735_index_offset_req_1 : boolean;
  signal array_obj_ref_1735_index_offset_ack_1 : boolean;
  signal phi_stmt_1828_req_1 : boolean;
  signal addr_of_1736_final_reg_req_0 : boolean;
  signal type_cast_1833_inst_ack_1 : boolean;
  signal addr_of_1736_final_reg_ack_0 : boolean;
  signal addr_of_1736_final_reg_req_1 : boolean;
  signal type_cast_1833_inst_req_1 : boolean;
  signal addr_of_1736_final_reg_ack_1 : boolean;
  signal type_cast_1831_inst_ack_0 : boolean;
  signal type_cast_1831_inst_req_0 : boolean;
  signal phi_stmt_1613_req_1 : boolean;
  signal type_cast_1619_inst_ack_1 : boolean;
  signal type_cast_1619_inst_req_1 : boolean;
  signal type_cast_1619_inst_ack_0 : boolean;
  signal type_cast_1833_inst_ack_0 : boolean;
  signal phi_stmt_1620_req_0 : boolean;
  signal type_cast_1619_inst_req_0 : boolean;
  signal type_cast_1833_inst_req_0 : boolean;
  signal ptr_deref_1739_store_0_req_0 : boolean;
  signal ptr_deref_1739_store_0_ack_0 : boolean;
  signal WPIPE_Block0_done_1844_inst_ack_1 : boolean;
  signal type_cast_1612_inst_ack_0 : boolean;
  signal ptr_deref_1739_store_0_req_1 : boolean;
  signal ptr_deref_1739_store_0_ack_1 : boolean;
  signal type_cast_1744_inst_req_0 : boolean;
  signal type_cast_1744_inst_ack_0 : boolean;
  signal type_cast_1744_inst_req_1 : boolean;
  signal type_cast_1744_inst_ack_1 : boolean;
  signal if_stmt_1757_branch_req_0 : boolean;
  signal if_stmt_1757_branch_ack_1 : boolean;
  signal if_stmt_1757_branch_ack_0 : boolean;
  signal type_cast_1785_inst_req_0 : boolean;
  signal type_cast_1785_inst_ack_0 : boolean;
  signal type_cast_1785_inst_req_1 : boolean;
  signal type_cast_1785_inst_ack_1 : boolean;
  signal type_cast_1801_inst_req_0 : boolean;
  signal type_cast_1801_inst_ack_0 : boolean;
  signal type_cast_1801_inst_req_1 : boolean;
  signal type_cast_1801_inst_ack_1 : boolean;
  signal if_stmt_1808_branch_req_0 : boolean;
  signal if_stmt_1808_branch_ack_1 : boolean;
  signal if_stmt_1808_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1844_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1844_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1844_inst_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3758_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3758_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3758_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3758_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3758: Block -- control-path 
    signal convTransposeA_CP_3758_elements: BooleanArray(125 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3758_elements(0) <= convTransposeA_CP_3758_start;
    convTransposeA_CP_3758_symbol <= convTransposeA_CP_3758_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1499_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1499_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1499_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1543_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1530_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/$entry
      -- CP-element group 0: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1543_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558__entry__
      -- CP-element group 0: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1543_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1497/branch_block_stmt_1497__entry__
      -- CP-element group 0: 	 branch_block_stmt_1497/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1530_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1530_update_start_
      -- 
    rr_3806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(0), ack => RPIPE_Block0_start_1499_inst_req_0); -- 
    cr_3979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(0), ack => type_cast_1543_inst_req_1); -- 
    cr_3951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(0), ack => type_cast_1530_inst_req_1); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	125 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	84 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	94 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1497/assign_stmt_1840__exit__
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_sources/type_cast_1619/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_sources/type_cast_1612/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1606/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/assign_stmt_1840__entry__
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_sources/type_cast_1612/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_sources/type_cast_1612/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/merge_stmt_1814__exit__
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_sources/type_cast_1612/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_sources/type_cast_1633/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_sources/type_cast_1633/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_sources/type_cast_1633/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_sources/type_cast_1633/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_sources/type_cast_1633/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_sources/type_cast_1633/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1627/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_sources/type_cast_1626/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_sources/type_cast_1626/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_sources/type_cast_1626/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1613/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_sources/type_cast_1612/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_sources/type_cast_1626/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_sources/type_cast_1626/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_sources/type_cast_1626/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1620/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_sources/type_cast_1619/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_sources/type_cast_1619/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_sources/type_cast_1619/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_sources/type_cast_1619/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_sources/type_cast_1612/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_sources/type_cast_1619/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/assign_stmt_1840/$entry
      -- CP-element group 1: 	 branch_block_stmt_1497/assign_stmt_1840/$exit
      -- 
    rr_4492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(1), ack => type_cast_1612_inst_req_0); -- 
    rr_4561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(1), ack => type_cast_1633_inst_req_0); -- 
    cr_4566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(1), ack => type_cast_1633_inst_req_1); -- 
    cr_4543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(1), ack => type_cast_1626_inst_req_1); -- 
    rr_4538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(1), ack => type_cast_1626_inst_req_0); -- 
    cr_4497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(1), ack => type_cast_1612_inst_req_1); -- 
    cr_4520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(1), ack => type_cast_1619_inst_req_1); -- 
    rr_4515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(1), ack => type_cast_1619_inst_req_0); -- 
    convTransposeA_CP_3758_elements(1) <= convTransposeA_CP_3758_elements(125);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1499_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1499_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1499_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1499_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1499_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1499_Update/cr
      -- 
    ra_3807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1499_inst_ack_0, ack => convTransposeA_CP_3758_elements(2)); -- 
    cr_3811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(2), ack => RPIPE_Block0_start_1499_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1502_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1499_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1499_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1502_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1499_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1502_sample_start_
      -- 
    ca_3812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1499_inst_ack_1, ack => convTransposeA_CP_3758_elements(3)); -- 
    rr_3820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(3), ack => RPIPE_Block0_start_1502_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1502_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1502_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1502_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1502_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1502_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1502_Sample/ra
      -- 
    ra_3821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1502_inst_ack_0, ack => convTransposeA_CP_3758_elements(4)); -- 
    cr_3825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(4), ack => RPIPE_Block0_start_1502_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1502_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1502_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1505_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1505_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1502_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1505_Sample/$entry
      -- 
    ca_3826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1502_inst_ack_1, ack => convTransposeA_CP_3758_elements(5)); -- 
    rr_3834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(5), ack => RPIPE_Block0_start_1505_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1505_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1505_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1505_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1505_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1505_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1505_Sample/$exit
      -- 
    ra_3835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1505_inst_ack_0, ack => convTransposeA_CP_3758_elements(6)); -- 
    cr_3839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(6), ack => RPIPE_Block0_start_1505_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1508_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1505_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1505_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1508_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1505_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1508_sample_start_
      -- 
    ca_3840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1505_inst_ack_1, ack => convTransposeA_CP_3758_elements(7)); -- 
    rr_3848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(7), ack => RPIPE_Block0_start_1508_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1508_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1508_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1508_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1508_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1508_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1508_Update/cr
      -- 
    ra_3849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1508_inst_ack_0, ack => convTransposeA_CP_3758_elements(8)); -- 
    cr_3853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(8), ack => RPIPE_Block0_start_1508_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1511_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1511_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1508_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1508_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1508_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1511_Sample/$entry
      -- 
    ca_3854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1508_inst_ack_1, ack => convTransposeA_CP_3758_elements(9)); -- 
    rr_3862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(9), ack => RPIPE_Block0_start_1511_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1511_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1511_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1511_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1511_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1511_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1511_Sample/$exit
      -- 
    ra_3863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1511_inst_ack_0, ack => convTransposeA_CP_3758_elements(10)); -- 
    cr_3867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(10), ack => RPIPE_Block0_start_1511_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1514_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1511_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1511_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1514_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1511_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1514_Sample/$entry
      -- 
    ca_3868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1511_inst_ack_1, ack => convTransposeA_CP_3758_elements(11)); -- 
    rr_3876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(11), ack => RPIPE_Block0_start_1514_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1514_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1514_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1514_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1514_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1514_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1514_Sample/$exit
      -- 
    ra_3877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1514_inst_ack_0, ack => convTransposeA_CP_3758_elements(12)); -- 
    cr_3881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(12), ack => RPIPE_Block0_start_1514_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1517_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1514_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1514_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1517_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1514_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1517_Sample/$entry
      -- 
    ca_3882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1514_inst_ack_1, ack => convTransposeA_CP_3758_elements(13)); -- 
    rr_3890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(13), ack => RPIPE_Block0_start_1517_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1517_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1517_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1517_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1517_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1517_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1517_update_start_
      -- 
    ra_3891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1517_inst_ack_0, ack => convTransposeA_CP_3758_elements(14)); -- 
    cr_3895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(14), ack => RPIPE_Block0_start_1517_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1517_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1517_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1520_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1517_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1520_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1520_Sample/rr
      -- 
    ca_3896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1517_inst_ack_1, ack => convTransposeA_CP_3758_elements(15)); -- 
    rr_3904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(15), ack => RPIPE_Block0_start_1520_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1520_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1520_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1520_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1520_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1520_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1520_Sample/ra
      -- 
    ra_3905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1520_inst_ack_0, ack => convTransposeA_CP_3758_elements(16)); -- 
    cr_3909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(16), ack => RPIPE_Block0_start_1520_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1523_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1520_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1523_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1520_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1520_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1523_Sample/$entry
      -- 
    ca_3910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1520_inst_ack_1, ack => convTransposeA_CP_3758_elements(17)); -- 
    rr_3918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(17), ack => RPIPE_Block0_start_1523_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1523_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1523_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1523_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1523_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1523_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1523_Update/cr
      -- 
    ra_3919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1523_inst_ack_0, ack => convTransposeA_CP_3758_elements(18)); -- 
    cr_3923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(18), ack => RPIPE_Block0_start_1523_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1523_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1526_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1523_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1523_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1526_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1526_Sample/rr
      -- 
    ca_3924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1523_inst_ack_1, ack => convTransposeA_CP_3758_elements(19)); -- 
    rr_3932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(19), ack => RPIPE_Block0_start_1526_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1526_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1526_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1526_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1526_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1526_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1526_Sample/ra
      -- 
    ra_3933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1526_inst_ack_0, ack => convTransposeA_CP_3758_elements(20)); -- 
    cr_3937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(20), ack => RPIPE_Block0_start_1526_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1530_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1530_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1539_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1539_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1539_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1526_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1530_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1526_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1526_Update/$exit
      -- 
    ca_3938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1526_inst_ack_1, ack => convTransposeA_CP_3758_elements(21)); -- 
    rr_3946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(21), ack => type_cast_1530_inst_req_0); -- 
    rr_3960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(21), ack => RPIPE_Block0_start_1539_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1530_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1530_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1530_sample_completed_
      -- 
    ra_3947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1530_inst_ack_0, ack => convTransposeA_CP_3758_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1530_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1530_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1530_Update/ca
      -- 
    ca_3952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1530_inst_ack_1, ack => convTransposeA_CP_3758_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1539_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1539_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1539_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1539_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1539_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1539_Sample/ra
      -- 
    ra_3961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1539_inst_ack_0, ack => convTransposeA_CP_3758_elements(24)); -- 
    cr_3965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(24), ack => RPIPE_Block0_start_1539_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1539_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1539_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1543_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1551_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1543_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1543_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1539_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1551_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1551_Sample/$entry
      -- 
    ca_3966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1539_inst_ack_1, ack => convTransposeA_CP_3758_elements(25)); -- 
    rr_3974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(25), ack => type_cast_1543_inst_req_0); -- 
    rr_3988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(25), ack => RPIPE_Block0_start_1551_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1543_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1543_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1543_Sample/ra
      -- 
    ra_3975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1543_inst_ack_0, ack => convTransposeA_CP_3758_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1543_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1543_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/type_cast_1543_Update/$exit
      -- 
    ca_3980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1543_inst_ack_1, ack => convTransposeA_CP_3758_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1551_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1551_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1551_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1551_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1551_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1551_Sample/$exit
      -- 
    ra_3989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1551_inst_ack_0, ack => convTransposeA_CP_3758_elements(28)); -- 
    cr_3993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(28), ack => RPIPE_Block0_start_1551_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1554_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1551_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1554_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1554_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1551_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1551_Update/$exit
      -- 
    ca_3994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1551_inst_ack_1, ack => convTransposeA_CP_3758_elements(29)); -- 
    rr_4002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(29), ack => RPIPE_Block0_start_1554_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1554_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1554_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1554_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1554_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1554_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1554_sample_completed_
      -- 
    ra_4003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1554_inst_ack_0, ack => convTransposeA_CP_3758_elements(30)); -- 
    cr_4007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(30), ack => RPIPE_Block0_start_1554_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1557_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1557_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1557_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1554_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1554_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1554_update_completed_
      -- 
    ca_4008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1554_inst_ack_1, ack => convTransposeA_CP_3758_elements(31)); -- 
    rr_4016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(31), ack => RPIPE_Block0_start_1557_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1557_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1557_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1557_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1557_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1557_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1557_Sample/$exit
      -- 
    ra_4017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1557_inst_ack_0, ack => convTransposeA_CP_3758_elements(32)); -- 
    cr_4021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(32), ack => RPIPE_Block0_start_1557_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1557_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1557_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/RPIPE_Block0_start_1557_Update/$exit
      -- 
    ca_4022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1557_inst_ack_1, ack => convTransposeA_CP_3758_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558__exit__
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1500_to_assign_stmt_1558/$exit
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603__entry__
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1592_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1592_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1588_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1592_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1592_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1588_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1588_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1588_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1588_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1588_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1584_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1584_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1584_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1584_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1584_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1584_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/$entry
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1592_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1592_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1596_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1596_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1596_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1596_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1596_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1596_Update/cr
      -- 
    cr_4052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(34), ack => type_cast_1588_inst_req_1); -- 
    rr_4061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(34), ack => type_cast_1592_inst_req_0); -- 
    rr_4047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(34), ack => type_cast_1588_inst_req_0); -- 
    cr_4038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(34), ack => type_cast_1584_inst_req_1); -- 
    rr_4033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(34), ack => type_cast_1584_inst_req_0); -- 
    cr_4066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(34), ack => type_cast_1592_inst_req_1); -- 
    rr_4075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(34), ack => type_cast_1596_inst_req_0); -- 
    cr_4080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(34), ack => type_cast_1596_inst_req_1); -- 
    convTransposeA_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(23) & convTransposeA_CP_3758_elements(27) & convTransposeA_CP_3758_elements(33);
      gj_convTransposeA_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1584_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1584_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1584_sample_completed_
      -- 
    ra_4034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1584_inst_ack_0, ack => convTransposeA_CP_3758_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1584_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1584_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1584_update_completed_
      -- 
    ca_4039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1584_inst_ack_1, ack => convTransposeA_CP_3758_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1588_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1588_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1588_sample_completed_
      -- 
    ra_4048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1588_inst_ack_0, ack => convTransposeA_CP_3758_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1588_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1588_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1588_update_completed_
      -- 
    ca_4053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1588_inst_ack_1, ack => convTransposeA_CP_3758_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1592_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1592_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1592_Sample/$exit
      -- 
    ra_4062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1592_inst_ack_0, ack => convTransposeA_CP_3758_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1592_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1592_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1592_Update/ca
      -- 
    ca_4067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1592_inst_ack_1, ack => convTransposeA_CP_3758_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1596_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1596_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1596_Sample/ra
      -- 
    ra_4076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1596_inst_ack_0, ack => convTransposeA_CP_3758_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1596_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1596_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/type_cast_1596_Update/ca
      -- 
    ca_4081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1596_inst_ack_1, ack => convTransposeA_CP_3758_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43:  members (12) 
      -- CP-element group 43: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603__exit__
      -- CP-element group 43: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1613/$entry
      -- CP-element group 43: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1497/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1620/$entry
      -- CP-element group 43: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1606/$entry
      -- CP-element group 43: 	 branch_block_stmt_1497/assign_stmt_1565_to_assign_stmt_1603/$exit
      -- CP-element group 43: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1627/$entry
      -- CP-element group 43: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/$entry
      -- 
    convTransposeA_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(36) & convTransposeA_CP_3758_elements(38) & convTransposeA_CP_3758_elements(40) & convTransposeA_CP_3758_elements(42);
      gj_convTransposeA_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	102 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1668_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1668_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1668_Sample/ra
      -- 
    ra_4093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1668_inst_ack_0, ack => convTransposeA_CP_3758_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	102 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1668_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1668_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1668_Update/ca
      -- 
    ca_4098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1668_inst_ack_1, ack => convTransposeA_CP_3758_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	102 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1672_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1672_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1672_Sample/ra
      -- 
    ra_4107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1672_inst_ack_0, ack => convTransposeA_CP_3758_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	102 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1672_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1672_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1672_Update/ca
      -- 
    ca_4112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1672_inst_ack_1, ack => convTransposeA_CP_3758_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	102 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1676_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1676_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1676_Sample/ra
      -- 
    ra_4121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1676_inst_ack_0, ack => convTransposeA_CP_3758_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	102 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1676_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1676_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1676_Update/ca
      -- 
    ca_4126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1676_inst_ack_1, ack => convTransposeA_CP_3758_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	102 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1706_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1706_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1706_Sample/ra
      -- 
    ra_4135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1706_inst_ack_0, ack => convTransposeA_CP_3758_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	102 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1706_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1706_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1706_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_final_index_sum_regn_Sample/req
      -- 
    ca_4140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1706_inst_ack_1, ack => convTransposeA_CP_3758_elements(51)); -- 
    req_4165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(51), ack => array_obj_ref_1712_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_final_index_sum_regn_Sample/ack
      -- 
    ack_4166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1712_index_offset_ack_0, ack => convTransposeA_CP_3758_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	102 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1713_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1713_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1713_request/req
      -- 
    ack_4171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1712_index_offset_ack_1, ack => convTransposeA_CP_3758_elements(53)); -- 
    req_4180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(53), ack => addr_of_1713_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1713_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1713_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1713_request/ack
      -- 
    ack_4181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1713_final_reg_ack_0, ack => convTransposeA_CP_3758_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	102 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1713_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1713_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1713_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Sample/word_access_start/word_0/rr
      -- 
    ack_4186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1713_final_reg_ack_1, ack => convTransposeA_CP_3758_elements(55)); -- 
    rr_4219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(55), ack => ptr_deref_1717_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Sample/word_access_start/word_0/ra
      -- 
    ra_4220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_load_0_ack_0, ack => convTransposeA_CP_3758_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	102 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Update/ptr_deref_1717_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Update/ptr_deref_1717_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Update/ptr_deref_1717_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Update/ptr_deref_1717_Merge/merge_ack
      -- 
    ca_4231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_load_0_ack_1, ack => convTransposeA_CP_3758_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_final_index_sum_regn_Sample/req
      -- 
    req_4261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(58), ack => array_obj_ref_1735_index_offset_req_0); -- 
    convTransposeA_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(45) & convTransposeA_CP_3758_elements(47) & convTransposeA_CP_3758_elements(49);
      gj_convTransposeA_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_final_index_sum_regn_Sample/ack
      -- 
    ack_4262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1735_index_offset_ack_0, ack => convTransposeA_CP_3758_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	102 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1736_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1736_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1736_request/req
      -- 
    ack_4267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1735_index_offset_ack_1, ack => convTransposeA_CP_3758_elements(60)); -- 
    req_4276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(60), ack => addr_of_1736_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1736_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1736_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1736_request/ack
      -- 
    ack_4277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1736_final_reg_ack_0, ack => convTransposeA_CP_3758_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	102 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1736_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1736_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1736_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_word_addrgen/root_register_ack
      -- 
    ack_4282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1736_final_reg_ack_1, ack => convTransposeA_CP_3758_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Sample/ptr_deref_1739_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Sample/ptr_deref_1739_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Sample/ptr_deref_1739_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Sample/ptr_deref_1739_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Sample/word_access_start/word_0/rr
      -- 
    rr_4320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(63), ack => ptr_deref_1739_store_0_req_0); -- 
    convTransposeA_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(57) & convTransposeA_CP_3758_elements(62);
      gj_convTransposeA_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Sample/word_access_start/word_0/ra
      -- 
    ra_4321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1739_store_0_ack_0, ack => convTransposeA_CP_3758_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	102 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Update/word_access_complete/word_0/ca
      -- 
    ca_4332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1739_store_0_ack_1, ack => convTransposeA_CP_3758_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	102 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1744_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1744_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1744_Sample/ra
      -- 
    ra_4341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1744_inst_ack_0, ack => convTransposeA_CP_3758_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	102 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1744_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1744_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1744_Update/ca
      -- 
    ca_4346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1744_inst_ack_1, ack => convTransposeA_CP_3758_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1497/if_stmt_1757__entry__
      -- CP-element group 68: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756__exit__
      -- CP-element group 68: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/$exit
      -- CP-element group 68: 	 branch_block_stmt_1497/if_stmt_1757_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1497/if_stmt_1757_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1497/if_stmt_1757_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1497/if_stmt_1757_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1497/R_cmp_1758_place
      -- CP-element group 68: 	 branch_block_stmt_1497/if_stmt_1757_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1497/if_stmt_1757_else_link/$entry
      -- 
    branch_req_4354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(68), ack => if_stmt_1757_branch_req_0); -- 
    convTransposeA_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(52) & convTransposeA_CP_3758_elements(59) & convTransposeA_CP_3758_elements(65) & convTransposeA_CP_3758_elements(67);
      gj_convTransposeA_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	111 
    -- CP-element group 69: 	112 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	115 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	118 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1497/merge_stmt_1763__exit__
      -- CP-element group 69: 	 branch_block_stmt_1497/assign_stmt_1769__entry__
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123
      -- CP-element group 69: 	 branch_block_stmt_1497/assign_stmt_1769__exit__
      -- CP-element group 69: 	 branch_block_stmt_1497/merge_stmt_1763_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1497/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1497/merge_stmt_1763_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1831/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1828/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1831/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_sources/type_cast_1821/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1831/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_sources/type_cast_1821/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/merge_stmt_1763_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_sources/type_cast_1821/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_sources/type_cast_1821/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_sources/type_cast_1821/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_sources/type_cast_1821/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/merge_stmt_1763_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1815/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1831/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1831/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1831/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1497/if_stmt_1757_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1497/if_stmt_1757_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1497/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1497/assign_stmt_1769/$entry
      -- CP-element group 69: 	 branch_block_stmt_1497/assign_stmt_1769/$exit
      -- 
    if_choice_transition_4359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1757_branch_ack_1, ack => convTransposeA_CP_3758_elements(69)); -- 
    cr_4727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(69), ack => type_cast_1821_inst_req_1); -- 
    rr_4722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(69), ack => type_cast_1821_inst_req_0); -- 
    cr_4704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(69), ack => type_cast_1827_inst_req_1); -- 
    rr_4699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(69), ack => type_cast_1827_inst_req_0); -- 
    cr_4681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(69), ack => type_cast_1831_inst_req_1); -- 
    rr_4676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(69), ack => type_cast_1831_inst_req_0); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1497/merge_stmt_1771__exit__
      -- CP-element group 70: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807__entry__
      -- CP-element group 70: 	 branch_block_stmt_1497/merge_stmt_1771_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1497/merge_stmt_1771_PhiAck/dummy
      -- CP-element group 70: 	 branch_block_stmt_1497/merge_stmt_1771_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1497/merge_stmt_1771_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1497/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1497/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1497/if_stmt_1757_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1497/if_stmt_1757_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1497/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/$entry
      -- CP-element group 70: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1785_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1785_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1785_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1785_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1785_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1785_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1801_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1801_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1801_Update/cr
      -- 
    else_choice_transition_4363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1757_branch_ack_0, ack => convTransposeA_CP_3758_elements(70)); -- 
    rr_4379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(70), ack => type_cast_1785_inst_req_0); -- 
    cr_4384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(70), ack => type_cast_1785_inst_req_1); -- 
    cr_4398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(70), ack => type_cast_1801_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1785_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1785_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1785_Sample/ra
      -- 
    ra_4380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1785_inst_ack_0, ack => convTransposeA_CP_3758_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1785_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1785_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1785_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1801_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1801_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1801_Sample/rr
      -- 
    ca_4385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1785_inst_ack_1, ack => convTransposeA_CP_3758_elements(72)); -- 
    rr_4393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(72), ack => type_cast_1801_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1801_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1801_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1801_Sample/ra
      -- 
    ra_4394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1801_inst_ack_0, ack => convTransposeA_CP_3758_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807__exit__
      -- CP-element group 74: 	 branch_block_stmt_1497/if_stmt_1808__entry__
      -- CP-element group 74: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/$exit
      -- CP-element group 74: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1801_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1801_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1497/assign_stmt_1777_to_assign_stmt_1807/type_cast_1801_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1497/if_stmt_1808_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1497/if_stmt_1808_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1497/if_stmt_1808_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1497/if_stmt_1808_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1497/R_cmp112_1809_place
      -- CP-element group 74: 	 branch_block_stmt_1497/if_stmt_1808_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1497/if_stmt_1808_else_link/$entry
      -- 
    ca_4399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1801_inst_ack_1, ack => convTransposeA_CP_3758_elements(74)); -- 
    branch_req_4407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(74), ack => if_stmt_1808_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1497/merge_stmt_1842__exit__
      -- CP-element group 75: 	 branch_block_stmt_1497/assign_stmt_1847__entry__
      -- CP-element group 75: 	 branch_block_stmt_1497/merge_stmt_1842_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1497/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1497/merge_stmt_1842_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1497/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1497/merge_stmt_1842_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_1497/merge_stmt_1842_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1497/if_stmt_1808_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1497/if_stmt_1808_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1497/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1497/assign_stmt_1847/$entry
      -- CP-element group 75: 	 branch_block_stmt_1497/assign_stmt_1847/WPIPE_Block0_done_1844_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1497/assign_stmt_1847/WPIPE_Block0_done_1844_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1497/assign_stmt_1847/WPIPE_Block0_done_1844_Sample/req
      -- 
    if_choice_transition_4412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1808_branch_ack_1, ack => convTransposeA_CP_3758_elements(75)); -- 
    req_4432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(75), ack => WPIPE_Block0_done_1844_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	103 
    -- CP-element group 76: 	104 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	109 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1833/$entry
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1828/$entry
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1833/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1833/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1815/$entry
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/$entry
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/$entry
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1833/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1833/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1833/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1497/if_stmt_1808_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1497/if_stmt_1808_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123
      -- 
    else_choice_transition_4416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1808_branch_ack_0, ack => convTransposeA_CP_3758_elements(76)); -- 
    cr_4647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(76), ack => type_cast_1825_inst_req_1); -- 
    rr_4642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(76), ack => type_cast_1825_inst_req_0); -- 
    cr_4624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(76), ack => type_cast_1833_inst_req_1); -- 
    rr_4619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(76), ack => type_cast_1833_inst_req_0); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1497/assign_stmt_1847/WPIPE_Block0_done_1844_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1497/assign_stmt_1847/WPIPE_Block0_done_1844_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1497/assign_stmt_1847/WPIPE_Block0_done_1844_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1497/assign_stmt_1847/WPIPE_Block0_done_1844_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1497/assign_stmt_1847/WPIPE_Block0_done_1844_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1497/assign_stmt_1847/WPIPE_Block0_done_1844_Update/req
      -- 
    ack_4433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1844_inst_ack_0, ack => convTransposeA_CP_3758_elements(77)); -- 
    req_4437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(77), ack => WPIPE_Block0_done_1844_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 branch_block_stmt_1497/merge_stmt_1849__exit__
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1497/branch_block_stmt_1497__exit__
      -- CP-element group 78: 	 branch_block_stmt_1497/$exit
      -- CP-element group 78: 	 branch_block_stmt_1497/return__
      -- CP-element group 78: 	 branch_block_stmt_1497/assign_stmt_1847__exit__
      -- CP-element group 78: 	 branch_block_stmt_1497/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1497/merge_stmt_1849_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1497/merge_stmt_1849_PhiAck/dummy
      -- CP-element group 78: 	 branch_block_stmt_1497/merge_stmt_1849_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1497/merge_stmt_1849_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1497/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1497/assign_stmt_1847/WPIPE_Block0_done_1844_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_1497/assign_stmt_1847/$exit
      -- CP-element group 78: 	 branch_block_stmt_1497/assign_stmt_1847/WPIPE_Block0_done_1844_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1497/assign_stmt_1847/WPIPE_Block0_done_1844_Update/$exit
      -- 
    ack_4438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1844_inst_ack_1, ack => convTransposeA_CP_3758_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	83 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1606/$exit
      -- CP-element group 79: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_sources/type_cast_1610_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_req
      -- CP-element group 79: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_sources/$exit
      -- 
    phi_stmt_1606_req_4449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1606_req_4449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(79), ack => phi_stmt_1606_req_0); -- 
    -- Element group convTransposeA_CP_3758_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeA_CP_3758_elements(43), ack => convTransposeA_CP_3758_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1613/$exit
      -- CP-element group 80: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_req
      -- CP-element group 80: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_sources/type_cast_1617_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_sources/$exit
      -- 
    phi_stmt_1613_req_4457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1613_req_4457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(80), ack => phi_stmt_1613_req_0); -- 
    -- Element group convTransposeA_CP_3758_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeA_CP_3758_elements(43), ack => convTransposeA_CP_3758_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  output  delay-element  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_sources/type_cast_1624_konst_delay_trans
      -- CP-element group 81: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1620/$exit
      -- CP-element group 81: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_req
      -- 
    phi_stmt_1620_req_4465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1620_req_4465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(81), ack => phi_stmt_1620_req_0); -- 
    -- Element group convTransposeA_CP_3758_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convTransposeA_CP_3758_elements(43), ack => convTransposeA_CP_3758_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_sources/type_cast_1631_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_req
      -- CP-element group 82: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/phi_stmt_1627/$exit
      -- 
    phi_stmt_1627_req_4473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1627_req_4473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(82), ack => phi_stmt_1627_req_0); -- 
    -- Element group convTransposeA_CP_3758_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeA_CP_3758_elements(43), ack => convTransposeA_CP_3758_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  join  transition  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	79 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	97 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1497/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(79) & convTransposeA_CP_3758_elements(80) & convTransposeA_CP_3758_elements(81) & convTransposeA_CP_3758_elements(82);
      gj_convTransposeA_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	1 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_sources/type_cast_1612/SplitProtocol/Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_sources/type_cast_1612/SplitProtocol/Sample/ra
      -- 
    ra_4493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1612_inst_ack_0, ack => convTransposeA_CP_3758_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_sources/type_cast_1612/SplitProtocol/Update/ca
      -- CP-element group 85: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_sources/type_cast_1612/SplitProtocol/Update/$exit
      -- 
    ca_4498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1612_inst_ack_1, ack => convTransposeA_CP_3758_elements(85)); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	96 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1606/$exit
      -- CP-element group 86: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_sources/type_cast_1612/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_sources/type_cast_1612/$exit
      -- CP-element group 86: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1606/phi_stmt_1606_req
      -- 
    phi_stmt_1606_req_4499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1606_req_4499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(86), ack => phi_stmt_1606_req_1); -- 
    convTransposeA_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(84) & convTransposeA_CP_3758_elements(85);
      gj_convTransposeA_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_sources/type_cast_1619/SplitProtocol/Sample/ra
      -- CP-element group 87: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_sources/type_cast_1619/SplitProtocol/Sample/$exit
      -- 
    ra_4516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1619_inst_ack_0, ack => convTransposeA_CP_3758_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_sources/type_cast_1619/SplitProtocol/Update/ca
      -- CP-element group 88: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_sources/type_cast_1619/SplitProtocol/Update/$exit
      -- 
    ca_4521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1619_inst_ack_1, ack => convTransposeA_CP_3758_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	96 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_sources/type_cast_1619/$exit
      -- CP-element group 89: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1613/$exit
      -- CP-element group 89: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_req
      -- CP-element group 89: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1613/phi_stmt_1613_sources/type_cast_1619/SplitProtocol/$exit
      -- 
    phi_stmt_1613_req_4522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1613_req_4522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(89), ack => phi_stmt_1613_req_1); -- 
    convTransposeA_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(87) & convTransposeA_CP_3758_elements(88);
      gj_convTransposeA_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_sources/type_cast_1626/SplitProtocol/Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_sources/type_cast_1626/SplitProtocol/Sample/$exit
      -- 
    ra_4539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1626_inst_ack_0, ack => convTransposeA_CP_3758_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_sources/type_cast_1626/SplitProtocol/Update/ca
      -- CP-element group 91: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_sources/type_cast_1626/SplitProtocol/Update/$exit
      -- 
    ca_4544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1626_inst_ack_1, ack => convTransposeA_CP_3758_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	96 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_req
      -- CP-element group 92: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_sources/type_cast_1626/SplitProtocol/$exit
      -- CP-element group 92: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_sources/type_cast_1626/$exit
      -- CP-element group 92: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1620/phi_stmt_1620_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1620/$exit
      -- 
    phi_stmt_1620_req_4545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1620_req_4545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(92), ack => phi_stmt_1620_req_1); -- 
    convTransposeA_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(90) & convTransposeA_CP_3758_elements(91);
      gj_convTransposeA_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_sources/type_cast_1633/SplitProtocol/Sample/ra
      -- CP-element group 93: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_sources/type_cast_1633/SplitProtocol/Sample/$exit
      -- 
    ra_4562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1633_inst_ack_0, ack => convTransposeA_CP_3758_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	1 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_sources/type_cast_1633/SplitProtocol/Update/ca
      -- CP-element group 94: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_sources/type_cast_1633/SplitProtocol/Update/$exit
      -- 
    ca_4567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1633_inst_ack_1, ack => convTransposeA_CP_3758_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_req
      -- CP-element group 95: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_sources/type_cast_1633/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_sources/type_cast_1633/$exit
      -- CP-element group 95: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1627/phi_stmt_1627_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/phi_stmt_1627/$exit
      -- 
    phi_stmt_1627_req_4568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1627_req_4568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(95), ack => phi_stmt_1627_req_1); -- 
    convTransposeA_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(93) & convTransposeA_CP_3758_elements(94);
      gj_convTransposeA_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	86 
    -- CP-element group 96: 	89 
    -- CP-element group 96: 	92 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_1497/ifx_xend123_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(86) & convTransposeA_CP_3758_elements(89) & convTransposeA_CP_3758_elements(92) & convTransposeA_CP_3758_elements(95);
      gj_convTransposeA_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  merge  fork  transition  place  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	83 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: 	99 
    -- CP-element group 97: 	100 
    -- CP-element group 97: 	101 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_1497/merge_stmt_1605_PhiAck/$entry
      -- CP-element group 97: 	 branch_block_stmt_1497/merge_stmt_1605_PhiReqMerge
      -- 
    convTransposeA_CP_3758_elements(97) <= OrReduce(convTransposeA_CP_3758_elements(83) & convTransposeA_CP_3758_elements(96));
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	102 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1497/merge_stmt_1605_PhiAck/phi_stmt_1606_ack
      -- 
    phi_stmt_1606_ack_4573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1606_ack_0, ack => convTransposeA_CP_3758_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1497/merge_stmt_1605_PhiAck/phi_stmt_1613_ack
      -- 
    phi_stmt_1613_ack_4574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1613_ack_0, ack => convTransposeA_CP_3758_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	97 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1497/merge_stmt_1605_PhiAck/phi_stmt_1620_ack
      -- 
    phi_stmt_1620_ack_4575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1620_ack_0, ack => convTransposeA_CP_3758_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	97 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1497/merge_stmt_1605_PhiAck/phi_stmt_1627_ack
      -- 
    phi_stmt_1627_ack_4576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1627_ack_0, ack => convTransposeA_CP_3758_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  place  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	98 
    -- CP-element group 102: 	99 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	44 
    -- CP-element group 102: 	45 
    -- CP-element group 102: 	46 
    -- CP-element group 102: 	47 
    -- CP-element group 102: 	48 
    -- CP-element group 102: 	49 
    -- CP-element group 102: 	50 
    -- CP-element group 102: 	51 
    -- CP-element group 102: 	53 
    -- CP-element group 102: 	55 
    -- CP-element group 102: 	57 
    -- CP-element group 102: 	60 
    -- CP-element group 102: 	62 
    -- CP-element group 102: 	65 
    -- CP-element group 102: 	66 
    -- CP-element group 102: 	67 
    -- CP-element group 102:  members (56) 
      -- CP-element group 102: 	 branch_block_stmt_1497/merge_stmt_1605_PhiAck/$exit
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756__entry__
      -- CP-element group 102: 	 branch_block_stmt_1497/merge_stmt_1605__exit__
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1668_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1668_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1668_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1668_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1668_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1668_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1672_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1672_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1672_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1672_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1672_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1672_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1676_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1676_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1676_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1676_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1676_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1676_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1706_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1706_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1706_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1706_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1706_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1706_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1713_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1712_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1713_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1713_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1717_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1736_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_final_index_sum_regn_update_start
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_final_index_sum_regn_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/array_obj_ref_1735_final_index_sum_regn_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1736_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/addr_of_1736_complete/req
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/ptr_deref_1739_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1744_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1744_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1744_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1744_Sample/rr
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1744_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1497/assign_stmt_1640_to_assign_stmt_1756/type_cast_1744_Update/cr
      -- 
    rr_4092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1668_inst_req_0); -- 
    cr_4097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1668_inst_req_1); -- 
    rr_4106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1672_inst_req_0); -- 
    cr_4111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1672_inst_req_1); -- 
    rr_4120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1676_inst_req_0); -- 
    cr_4125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1676_inst_req_1); -- 
    rr_4134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1706_inst_req_0); -- 
    cr_4139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1706_inst_req_1); -- 
    req_4170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => array_obj_ref_1712_index_offset_req_1); -- 
    req_4185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => addr_of_1713_final_reg_req_1); -- 
    cr_4230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => ptr_deref_1717_load_0_req_1); -- 
    req_4266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => array_obj_ref_1735_index_offset_req_1); -- 
    req_4281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => addr_of_1736_final_reg_req_1); -- 
    cr_4331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => ptr_deref_1739_store_0_req_1); -- 
    rr_4340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1744_inst_req_0); -- 
    cr_4345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(102), ack => type_cast_1744_inst_req_1); -- 
    convTransposeA_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(98) & convTransposeA_CP_3758_elements(99) & convTransposeA_CP_3758_elements(100) & convTransposeA_CP_3758_elements(101);
      gj_convTransposeA_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	76 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1833/SplitProtocol/Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1833/SplitProtocol/Sample/$exit
      -- 
    ra_4620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1833_inst_ack_0, ack => convTransposeA_CP_3758_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	76 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1833/SplitProtocol/Update/ca
      -- CP-element group 104: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1833/SplitProtocol/Update/$exit
      -- 
    ca_4625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1833_inst_ack_1, ack => convTransposeA_CP_3758_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	110 
    -- CP-element group 105:  members (5) 
      -- CP-element group 105: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1833/$exit
      -- CP-element group 105: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1833/SplitProtocol/$exit
      -- CP-element group 105: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1828/$exit
      -- CP-element group 105: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_req
      -- 
    phi_stmt_1828_req_4626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1828_req_4626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(105), ack => phi_stmt_1828_req_1); -- 
    convTransposeA_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(103) & convTransposeA_CP_3758_elements(104);
      gj_convTransposeA_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/Sample/$exit
      -- 
    ra_4643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1825_inst_ack_0, ack => convTransposeA_CP_3758_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/Update/ca
      -- CP-element group 107: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/Update/$exit
      -- 
    ca_4648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1825_inst_ack_1, ack => convTransposeA_CP_3758_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_req
      -- CP-element group 108: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1825/$exit
      -- CP-element group 108: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1822/$exit
      -- 
    phi_stmt_1822_req_4649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1822_req_4649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(108), ack => phi_stmt_1822_req_0); -- 
    convTransposeA_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(106) & convTransposeA_CP_3758_elements(107);
      gj_convTransposeA_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  output  delay-element  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_req
      -- CP-element group 109: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_sources/type_cast_1819_konst_delay_trans
      -- CP-element group 109: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_sources/$exit
      -- CP-element group 109: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/phi_stmt_1815/$exit
      -- 
    phi_stmt_1815_req_4657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1815_req_4657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(109), ack => phi_stmt_1815_req_0); -- 
    -- Element group convTransposeA_CP_3758_elements(109) is a control-delay.
    cp_element_109_delay: control_delay_element  generic map(name => " 109_delay", delay_value => 1)  port map(req => convTransposeA_CP_3758_elements(76), ack => convTransposeA_CP_3758_elements(109), clk => clk, reset =>reset);
    -- CP-element group 110:  join  transition  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	105 
    -- CP-element group 110: 	108 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	121 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1497/ifx_xelse_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(105) & convTransposeA_CP_3758_elements(108) & convTransposeA_CP_3758_elements(109);
      gj_convTransposeA_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	69 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1831/SplitProtocol/Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1831/SplitProtocol/Sample/$exit
      -- 
    ra_4677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1831_inst_ack_0, ack => convTransposeA_CP_3758_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	69 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1831/SplitProtocol/Update/ca
      -- CP-element group 112: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1831/SplitProtocol/Update/$exit
      -- 
    ca_4682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1831_inst_ack_1, ack => convTransposeA_CP_3758_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	120 
    -- CP-element group 113:  members (5) 
      -- CP-element group 113: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1831/$exit
      -- CP-element group 113: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/type_cast_1831/SplitProtocol/$exit
      -- CP-element group 113: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_sources/$exit
      -- CP-element group 113: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1828/$exit
      -- CP-element group 113: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1828/phi_stmt_1828_req
      -- 
    phi_stmt_1828_req_4683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1828_req_4683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(113), ack => phi_stmt_1828_req_0); -- 
    convTransposeA_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(111) & convTransposeA_CP_3758_elements(112);
      gj_convTransposeA_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/Sample/$exit
      -- 
    ra_4700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1827_inst_ack_0, ack => convTransposeA_CP_3758_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	69 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/Update/ca
      -- CP-element group 115: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/Update/$exit
      -- 
    ca_4705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1827_inst_ack_1, ack => convTransposeA_CP_3758_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	120 
    -- CP-element group 116:  members (5) 
      -- CP-element group 116: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_req
      -- CP-element group 116: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/SplitProtocol/$exit
      -- CP-element group 116: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/type_cast_1827/$exit
      -- CP-element group 116: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/phi_stmt_1822_sources/$exit
      -- CP-element group 116: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1822/$exit
      -- 
    phi_stmt_1822_req_4706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1822_req_4706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(116), ack => phi_stmt_1822_req_1); -- 
    convTransposeA_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(114) & convTransposeA_CP_3758_elements(115);
      gj_convTransposeA_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_sources/type_cast_1821/SplitProtocol/Sample/ra
      -- CP-element group 117: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_sources/type_cast_1821/SplitProtocol/Sample/$exit
      -- 
    ra_4723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1821_inst_ack_0, ack => convTransposeA_CP_3758_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	69 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_sources/type_cast_1821/SplitProtocol/Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_sources/type_cast_1821/SplitProtocol/Update/ca
      -- 
    ca_4728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1821_inst_ack_1, ack => convTransposeA_CP_3758_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_req
      -- CP-element group 119: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_sources/type_cast_1821/SplitProtocol/$exit
      -- CP-element group 119: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_sources/type_cast_1821/$exit
      -- CP-element group 119: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1815/phi_stmt_1815_sources/$exit
      -- CP-element group 119: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/phi_stmt_1815/$exit
      -- 
    phi_stmt_1815_req_4729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1815_req_4729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3758_elements(119), ack => phi_stmt_1815_req_1); -- 
    convTransposeA_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(117) & convTransposeA_CP_3758_elements(118);
      gj_convTransposeA_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	113 
    -- CP-element group 120: 	116 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_1497/ifx_xthen_ifx_xend123_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(113) & convTransposeA_CP_3758_elements(116) & convTransposeA_CP_3758_elements(119);
      gj_convTransposeA_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  merge  fork  transition  place  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	110 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: 	123 
    -- CP-element group 121: 	124 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_1497/merge_stmt_1814_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_1497/merge_stmt_1814_PhiReqMerge
      -- 
    convTransposeA_CP_3758_elements(121) <= OrReduce(convTransposeA_CP_3758_elements(110) & convTransposeA_CP_3758_elements(120));
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	125 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1497/merge_stmt_1814_PhiAck/phi_stmt_1815_ack
      -- 
    phi_stmt_1815_ack_4734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1815_ack_0, ack => convTransposeA_CP_3758_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1497/merge_stmt_1814_PhiAck/phi_stmt_1822_ack
      -- 
    phi_stmt_1822_ack_4735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1822_ack_0, ack => convTransposeA_CP_3758_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1497/merge_stmt_1814_PhiAck/phi_stmt_1828_ack
      -- 
    phi_stmt_1828_ack_4736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1828_ack_0, ack => convTransposeA_CP_3758_elements(124)); -- 
    -- CP-element group 125:  join  transition  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	122 
    -- CP-element group 125: 	123 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	1 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1497/merge_stmt_1814_PhiAck/$exit
      -- 
    convTransposeA_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3758_elements(122) & convTransposeA_CP_3758_elements(123) & convTransposeA_CP_3758_elements(124);
      gj_convTransposeA_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3758_elements(125), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom81_1734_resized : std_logic_vector(13 downto 0);
    signal R_idxprom81_1734_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1711_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1711_scaled : std_logic_vector(13 downto 0);
    signal add41_1565 : std_logic_vector(15 downto 0);
    signal add54_1576 : std_logic_vector(15 downto 0);
    signal add73_1687 : std_logic_vector(63 downto 0);
    signal add75_1697 : std_logic_vector(63 downto 0);
    signal add86_1751 : std_logic_vector(31 downto 0);
    signal add93_1769 : std_logic_vector(15 downto 0);
    signal add_1549 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_1645 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1712_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1712_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1712_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1712_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1712_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1712_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1735_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1735_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1735_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1735_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1735_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1735_root_address : std_logic_vector(13 downto 0);
    signal arrayidx77_1714 : std_logic_vector(31 downto 0);
    signal arrayidx82_1737 : std_logic_vector(31 downto 0);
    signal call11_1518 : std_logic_vector(15 downto 0);
    signal call13_1521 : std_logic_vector(15 downto 0);
    signal call14_1524 : std_logic_vector(15 downto 0);
    signal call15_1527 : std_logic_vector(15 downto 0);
    signal call16_1540 : std_logic_vector(15 downto 0);
    signal call18_1552 : std_logic_vector(15 downto 0);
    signal call1_1503 : std_logic_vector(15 downto 0);
    signal call20_1555 : std_logic_vector(15 downto 0);
    signal call22_1558 : std_logic_vector(15 downto 0);
    signal call3_1506 : std_logic_vector(15 downto 0);
    signal call5_1509 : std_logic_vector(15 downto 0);
    signal call7_1512 : std_logic_vector(15 downto 0);
    signal call9_1515 : std_logic_vector(15 downto 0);
    signal call_1500 : std_logic_vector(15 downto 0);
    signal cmp101_1782 : std_logic_vector(0 downto 0);
    signal cmp112_1807 : std_logic_vector(0 downto 0);
    signal cmp_1756 : std_logic_vector(0 downto 0);
    signal conv107_1802 : std_logic_vector(31 downto 0);
    signal conv110_1597 : std_logic_vector(31 downto 0);
    signal conv17_1544 : std_logic_vector(31 downto 0);
    signal conv61_1669 : std_logic_vector(63 downto 0);
    signal conv64_1585 : std_logic_vector(63 downto 0);
    signal conv66_1673 : std_logic_vector(63 downto 0);
    signal conv69_1589 : std_logic_vector(63 downto 0);
    signal conv71_1677 : std_logic_vector(63 downto 0);
    signal conv85_1745 : std_logic_vector(31 downto 0);
    signal conv89_1593 : std_logic_vector(31 downto 0);
    signal conv_1531 : std_logic_vector(31 downto 0);
    signal idxprom81_1730 : std_logic_vector(63 downto 0);
    signal idxprom_1707 : std_logic_vector(63 downto 0);
    signal inc105_1786 : std_logic_vector(15 downto 0);
    signal inc105x_xinput_dim0x_x2_1791 : std_logic_vector(15 downto 0);
    signal inc_1777 : std_logic_vector(15 downto 0);
    signal indvar_1606 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_1840 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_1828 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1627 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_1822 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1620 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1798 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_1815 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1613 : std_logic_vector(15 downto 0);
    signal mul50_1660 : std_logic_vector(15 downto 0);
    signal mul72_1682 : std_logic_vector(63 downto 0);
    signal mul74_1692 : std_logic_vector(63 downto 0);
    signal mul_1650 : std_logic_vector(15 downto 0);
    signal ptr_deref_1717_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1717_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1717_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1717_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1717_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1739_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1739_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1739_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1739_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1739_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1739_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1537 : std_logic_vector(31 downto 0);
    signal shr111126_1603 : std_logic_vector(31 downto 0);
    signal shr80_1724 : std_logic_vector(63 downto 0);
    signal shr_1703 : std_logic_vector(31 downto 0);
    signal sub44_1655 : std_logic_vector(15 downto 0);
    signal sub57_1581 : std_logic_vector(15 downto 0);
    signal sub58_1665 : std_logic_vector(15 downto 0);
    signal sub_1570 : std_logic_vector(15 downto 0);
    signal tmp1_1640 : std_logic_vector(31 downto 0);
    signal tmp78_1718 : std_logic_vector(63 downto 0);
    signal type_cast_1535_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1563_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1574_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1601_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1610_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1612_wire : std_logic_vector(31 downto 0);
    signal type_cast_1617_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1619_wire : std_logic_vector(15 downto 0);
    signal type_cast_1624_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1626_wire : std_logic_vector(15 downto 0);
    signal type_cast_1631_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1633_wire : std_logic_vector(15 downto 0);
    signal type_cast_1638_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1701_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1722_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1728_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1749_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1767_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1775_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1795_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1819_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1821_wire : std_logic_vector(15 downto 0);
    signal type_cast_1825_wire : std_logic_vector(15 downto 0);
    signal type_cast_1827_wire : std_logic_vector(15 downto 0);
    signal type_cast_1831_wire : std_logic_vector(15 downto 0);
    signal type_cast_1833_wire : std_logic_vector(15 downto 0);
    signal type_cast_1838_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1846_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_1712_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1712_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1712_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1712_resized_base_address <= "00000000000000";
    array_obj_ref_1735_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1735_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1735_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1735_resized_base_address <= "00000000000000";
    ptr_deref_1717_word_offset_0 <= "00000000000000";
    ptr_deref_1739_word_offset_0 <= "00000000000000";
    type_cast_1535_wire_constant <= "00000000000000000000000000010000";
    type_cast_1563_wire_constant <= "1111111111111111";
    type_cast_1574_wire_constant <= "1111111111111111";
    type_cast_1601_wire_constant <= "00000000000000000000000000000010";
    type_cast_1610_wire_constant <= "00000000000000000000000000000000";
    type_cast_1617_wire_constant <= "0000000000000000";
    type_cast_1624_wire_constant <= "0000000000000000";
    type_cast_1631_wire_constant <= "0000000000000000";
    type_cast_1638_wire_constant <= "00000000000000000000000000000100";
    type_cast_1701_wire_constant <= "00000000000000000000000000000010";
    type_cast_1722_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1728_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_1749_wire_constant <= "00000000000000000000000000000100";
    type_cast_1767_wire_constant <= "0000000000000100";
    type_cast_1775_wire_constant <= "0000000000000001";
    type_cast_1795_wire_constant <= "0000000000000000";
    type_cast_1819_wire_constant <= "0000000000000000";
    type_cast_1838_wire_constant <= "00000000000000000000000000000001";
    type_cast_1846_wire_constant <= "0000000000000001";
    phi_stmt_1606: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1610_wire_constant & type_cast_1612_wire;
      req <= phi_stmt_1606_req_0 & phi_stmt_1606_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1606",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1606_ack_0,
          idata => idata,
          odata => indvar_1606,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1606
    phi_stmt_1613: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1617_wire_constant & type_cast_1619_wire;
      req <= phi_stmt_1613_req_0 & phi_stmt_1613_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1613",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1613_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1613,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1613
    phi_stmt_1620: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1624_wire_constant & type_cast_1626_wire;
      req <= phi_stmt_1620_req_0 & phi_stmt_1620_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1620",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1620_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1620,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1620
    phi_stmt_1627: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1631_wire_constant & type_cast_1633_wire;
      req <= phi_stmt_1627_req_0 & phi_stmt_1627_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1627",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1627_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1627,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1627
    phi_stmt_1815: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1819_wire_constant & type_cast_1821_wire;
      req <= phi_stmt_1815_req_0 & phi_stmt_1815_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1815",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1815_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_1815,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1815
    phi_stmt_1822: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1825_wire & type_cast_1827_wire;
      req <= phi_stmt_1822_req_0 & phi_stmt_1822_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1822",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1822_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_1822,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1822
    phi_stmt_1828: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1831_wire & type_cast_1833_wire;
      req <= phi_stmt_1828_req_0 & phi_stmt_1828_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1828",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1828_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_1828,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1828
    -- flow-through select operator MUX_1797_inst
    input_dim1x_x2_1798 <= type_cast_1795_wire_constant when (cmp101_1782(0) /=  '0') else inc_1777;
    addr_of_1713_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1713_final_reg_req_0;
      addr_of_1713_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1713_final_reg_req_1;
      addr_of_1713_final_reg_ack_1<= rack(0);
      addr_of_1713_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1713_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1712_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx77_1714,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1736_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1736_final_reg_req_0;
      addr_of_1736_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1736_final_reg_req_1;
      addr_of_1736_final_reg_ack_1<= rack(0);
      addr_of_1736_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1736_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1735_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_1737,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1530_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1530_inst_req_0;
      type_cast_1530_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1530_inst_req_1;
      type_cast_1530_inst_ack_1<= rack(0);
      type_cast_1530_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1530_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1527,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1531,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1543_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1543_inst_req_0;
      type_cast_1543_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1543_inst_req_1;
      type_cast_1543_inst_ack_1<= rack(0);
      type_cast_1543_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1543_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1540,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1544,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1584_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1584_inst_req_0;
      type_cast_1584_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1584_inst_req_1;
      type_cast_1584_inst_ack_1<= rack(0);
      type_cast_1584_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1584_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1558,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_1585,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1588_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1588_inst_req_0;
      type_cast_1588_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1588_inst_req_1;
      type_cast_1588_inst_ack_1<= rack(0);
      type_cast_1588_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1588_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1555,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_1589,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1592_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1592_inst_req_0;
      type_cast_1592_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1592_inst_req_1;
      type_cast_1592_inst_ack_1<= rack(0);
      type_cast_1592_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1592_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1506,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv89_1593,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1596_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1596_inst_req_0;
      type_cast_1596_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1596_inst_req_1;
      type_cast_1596_inst_ack_1<= rack(0);
      type_cast_1596_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1596_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1500,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_1597,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1612_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1612_inst_req_0;
      type_cast_1612_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1612_inst_req_1;
      type_cast_1612_inst_ack_1<= rack(0);
      type_cast_1612_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1612_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1840,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1612_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1619_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1619_inst_req_0;
      type_cast_1619_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1619_inst_req_1;
      type_cast_1619_inst_ack_1<= rack(0);
      type_cast_1619_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1619_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_1815,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1619_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1626_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1626_inst_req_0;
      type_cast_1626_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1626_inst_req_1;
      type_cast_1626_inst_ack_1<= rack(0);
      type_cast_1626_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1626_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_1822,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1626_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1633_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1633_inst_req_0;
      type_cast_1633_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1633_inst_req_1;
      type_cast_1633_inst_ack_1<= rack(0);
      type_cast_1633_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1633_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_1828,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1633_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1668_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1668_inst_req_0;
      type_cast_1668_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1668_inst_req_1;
      type_cast_1668_inst_ack_1<= rack(0);
      type_cast_1668_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1668_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1613,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_1669,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1672_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1672_inst_req_0;
      type_cast_1672_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1672_inst_req_1;
      type_cast_1672_inst_ack_1<= rack(0);
      type_cast_1672_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1672_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub58_1665,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1673,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1676_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1676_inst_req_0;
      type_cast_1676_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1676_inst_req_1;
      type_cast_1676_inst_ack_1<= rack(0);
      type_cast_1676_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1676_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub44_1655,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_1677,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1706_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1706_inst_req_0;
      type_cast_1706_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1706_inst_req_1;
      type_cast_1706_inst_ack_1<= rack(0);
      type_cast_1706_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1706_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_1703,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1707,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1744_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1744_inst_req_0;
      type_cast_1744_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1744_inst_req_1;
      type_cast_1744_inst_ack_1<= rack(0);
      type_cast_1744_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1744_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1613,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_1745,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1785_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1785_inst_req_0;
      type_cast_1785_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1785_inst_req_1;
      type_cast_1785_inst_ack_1<= rack(0);
      type_cast_1785_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1785_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp101_1782,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc105_1786,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1801_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1801_inst_req_0;
      type_cast_1801_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1801_inst_req_1;
      type_cast_1801_inst_ack_1<= rack(0);
      type_cast_1801_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1801_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1791,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_1802,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1821_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1821_inst_req_0;
      type_cast_1821_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1821_inst_req_1;
      type_cast_1821_inst_ack_1<= rack(0);
      type_cast_1821_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1821_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add93_1769,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1821_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1825_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1825_inst_req_0;
      type_cast_1825_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1825_inst_req_1;
      type_cast_1825_inst_ack_1<= rack(0);
      type_cast_1825_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1825_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1798,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1825_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1827_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1827_inst_req_0;
      type_cast_1827_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1827_inst_req_1;
      type_cast_1827_inst_ack_1<= rack(0);
      type_cast_1827_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1827_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1620,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1827_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1831_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1831_inst_req_0;
      type_cast_1831_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1831_inst_req_1;
      type_cast_1831_inst_ack_1<= rack(0);
      type_cast_1831_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1831_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1627,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1831_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1833_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1833_inst_req_0;
      type_cast_1833_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1833_inst_req_1;
      type_cast_1833_inst_ack_1<= rack(0);
      type_cast_1833_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1833_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc105x_xinput_dim0x_x2_1791,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1833_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1712_index_1_rename
    process(R_idxprom_1711_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1711_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1711_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1712_index_1_resize
    process(idxprom_1707) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1707;
      ov := iv(13 downto 0);
      R_idxprom_1711_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1712_root_address_inst
    process(array_obj_ref_1712_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1712_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1712_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1735_index_1_rename
    process(R_idxprom81_1734_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom81_1734_resized;
      ov(13 downto 0) := iv;
      R_idxprom81_1734_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1735_index_1_resize
    process(idxprom81_1730) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom81_1730;
      ov := iv(13 downto 0);
      R_idxprom81_1734_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1735_root_address_inst
    process(array_obj_ref_1735_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1735_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1735_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1717_addr_0
    process(ptr_deref_1717_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1717_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1717_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1717_base_resize
    process(arrayidx77_1714) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx77_1714;
      ov := iv(13 downto 0);
      ptr_deref_1717_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1717_gather_scatter
    process(ptr_deref_1717_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1717_data_0;
      ov(63 downto 0) := iv;
      tmp78_1718 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1717_root_address_inst
    process(ptr_deref_1717_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1717_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1717_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1739_addr_0
    process(ptr_deref_1739_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1739_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1739_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1739_base_resize
    process(arrayidx82_1737) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_1737;
      ov := iv(13 downto 0);
      ptr_deref_1739_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1739_gather_scatter
    process(tmp78_1718) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp78_1718;
      ov(63 downto 0) := iv;
      ptr_deref_1739_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1739_root_address_inst
    process(ptr_deref_1739_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1739_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1739_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1757_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1756;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1757_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1757_branch_req_0,
          ack0 => if_stmt_1757_branch_ack_0,
          ack1 => if_stmt_1757_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1808_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp112_1807;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1808_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1808_branch_req_0,
          ack0 => if_stmt_1808_branch_ack_0,
          ack1 => if_stmt_1808_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1564_inst
    process(call7_1512) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1512, type_cast_1563_wire_constant, tmp_var);
      add41_1565 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1575_inst
    process(call9_1515) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1515, type_cast_1574_wire_constant, tmp_var);
      add54_1576 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1654_inst
    process(sub_1570, mul_1650) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1570, mul_1650, tmp_var);
      sub44_1655 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1664_inst
    process(sub57_1581, mul50_1660) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub57_1581, mul50_1660, tmp_var);
      sub58_1665 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1768_inst
    process(input_dim2x_x1_1613) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1613, type_cast_1767_wire_constant, tmp_var);
      add93_1769 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1776_inst
    process(input_dim1x_x1_1620) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1620, type_cast_1775_wire_constant, tmp_var);
      inc_1777 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1790_inst
    process(inc105_1786, input_dim0x_x2_1627) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc105_1786, input_dim0x_x2_1627, tmp_var);
      inc105x_xinput_dim0x_x2_1791 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1644_inst
    process(add_1549, tmp1_1640) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1549, tmp1_1640, tmp_var);
      add_src_0x_x0_1645 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1750_inst
    process(conv85_1745) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv85_1745, type_cast_1749_wire_constant, tmp_var);
      add86_1751 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1839_inst
    process(indvar_1606) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1606, type_cast_1838_wire_constant, tmp_var);
      indvarx_xnext_1840 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1686_inst
    process(mul72_1682, conv66_1673) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul72_1682, conv66_1673, tmp_var);
      add73_1687 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1696_inst
    process(mul74_1692, conv61_1669) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul74_1692, conv61_1669, tmp_var);
      add75_1697 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1729_inst
    process(shr80_1724) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr80_1724, type_cast_1728_wire_constant, tmp_var);
      idxprom81_1730 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1781_inst
    process(inc_1777, call1_1503) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_1777, call1_1503, tmp_var);
      cmp101_1782 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1806_inst
    process(conv107_1802, shr111126_1603) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv107_1802, shr111126_1603, tmp_var);
      cmp112_1807 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1602_inst
    process(conv110_1597) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv110_1597, type_cast_1601_wire_constant, tmp_var);
      shr111126_1603 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1702_inst
    process(add_src_0x_x0_1645) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_1645, type_cast_1701_wire_constant, tmp_var);
      shr_1703 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1723_inst
    process(add75_1697) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add75_1697, type_cast_1722_wire_constant, tmp_var);
      shr80_1724 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1649_inst
    process(input_dim0x_x2_1627, call13_1521) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1627, call13_1521, tmp_var);
      mul_1650 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1659_inst
    process(input_dim1x_x1_1620, call13_1521) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1620, call13_1521, tmp_var);
      mul50_1660 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1639_inst
    process(indvar_1606) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1606, type_cast_1638_wire_constant, tmp_var);
      tmp1_1640 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1681_inst
    process(conv71_1677, conv69_1589) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv71_1677, conv69_1589, tmp_var);
      mul72_1682 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1691_inst
    process(add73_1687, conv64_1585) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_1687, conv64_1585, tmp_var);
      mul74_1692 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1548_inst
    process(shl_1537, conv17_1544) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1537, conv17_1544, tmp_var);
      add_1549 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1536_inst
    process(conv_1531) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1531, type_cast_1535_wire_constant, tmp_var);
      shl_1537 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1569_inst
    process(add41_1565, call14_1524) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add41_1565, call14_1524, tmp_var);
      sub_1570 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1580_inst
    process(add54_1576, call14_1524) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add54_1576, call14_1524, tmp_var);
      sub57_1581 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1755_inst
    process(add86_1751, conv89_1593) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add86_1751, conv89_1593, tmp_var);
      cmp_1756 <= tmp_var; --
    end process;
    -- shared split operator group (28) : array_obj_ref_1712_index_offset 
    ApIntAdd_group_28: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1711_scaled;
      array_obj_ref_1712_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1712_index_offset_req_0;
      array_obj_ref_1712_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1712_index_offset_req_1;
      array_obj_ref_1712_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_28_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : array_obj_ref_1735_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom81_1734_scaled;
      array_obj_ref_1735_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1735_index_offset_req_0;
      array_obj_ref_1735_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1735_index_offset_req_1;
      array_obj_ref_1735_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared load operator group (0) : ptr_deref_1717_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1717_load_0_req_0;
      ptr_deref_1717_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1717_load_0_req_1;
      ptr_deref_1717_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1717_word_address_0;
      ptr_deref_1717_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1739_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1739_store_0_req_0;
      ptr_deref_1739_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1739_store_0_req_1;
      ptr_deref_1739_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1739_word_address_0;
      data_in <= ptr_deref_1739_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1511_inst RPIPE_Block0_start_1523_inst RPIPE_Block0_start_1539_inst RPIPE_Block0_start_1505_inst RPIPE_Block0_start_1520_inst RPIPE_Block0_start_1517_inst RPIPE_Block0_start_1514_inst RPIPE_Block0_start_1502_inst RPIPE_Block0_start_1508_inst RPIPE_Block0_start_1551_inst RPIPE_Block0_start_1499_inst RPIPE_Block0_start_1526_inst RPIPE_Block0_start_1557_inst RPIPE_Block0_start_1554_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block0_start_1511_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block0_start_1523_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block0_start_1539_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block0_start_1505_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block0_start_1520_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block0_start_1517_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block0_start_1514_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block0_start_1502_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_start_1508_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_start_1551_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_start_1499_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_start_1526_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_start_1557_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_start_1554_inst_req_0;
      RPIPE_Block0_start_1511_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block0_start_1523_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block0_start_1539_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block0_start_1505_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block0_start_1520_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block0_start_1517_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block0_start_1514_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block0_start_1502_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_start_1508_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_start_1551_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_start_1499_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_start_1526_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_start_1557_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_start_1554_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block0_start_1511_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block0_start_1523_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block0_start_1539_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block0_start_1505_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block0_start_1520_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block0_start_1517_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block0_start_1514_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block0_start_1502_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_start_1508_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_start_1551_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_start_1499_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_start_1526_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_start_1557_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_start_1554_inst_req_1;
      RPIPE_Block0_start_1511_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block0_start_1523_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block0_start_1539_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block0_start_1505_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block0_start_1520_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block0_start_1517_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block0_start_1514_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block0_start_1502_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_start_1508_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_start_1551_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_start_1499_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_start_1526_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_start_1557_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_start_1554_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call7_1512 <= data_out(223 downto 208);
      call14_1524 <= data_out(207 downto 192);
      call16_1540 <= data_out(191 downto 176);
      call3_1506 <= data_out(175 downto 160);
      call13_1521 <= data_out(159 downto 144);
      call11_1518 <= data_out(143 downto 128);
      call9_1515 <= data_out(127 downto 112);
      call1_1503 <= data_out(111 downto 96);
      call5_1509 <= data_out(95 downto 80);
      call18_1552 <= data_out(79 downto 64);
      call_1500 <= data_out(63 downto 48);
      call15_1527 <= data_out(47 downto 32);
      call22_1558 <= data_out(31 downto 16);
      call20_1555 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1844_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1844_inst_req_0;
      WPIPE_Block0_done_1844_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1844_inst_req_1;
      WPIPE_Block0_done_1844_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1846_wire_constant;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_4753_start: Boolean;
  signal convTransposeB_CP_4753_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block1_start_1870_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1870_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1895_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1864_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1858_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1895_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1870_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1858_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1870_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1867_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1873_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1864_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1867_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1858_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1864_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1910_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1910_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1910_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1907_inst_req_1 : boolean;
  signal type_cast_1899_inst_req_0 : boolean;
  signal type_cast_1899_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1879_inst_ack_1 : boolean;
  signal phi_stmt_2189_req_1 : boolean;
  signal RPIPE_Block1_start_1913_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1913_inst_ack_1 : boolean;
  signal type_cast_2194_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1895_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1907_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1907_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1879_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1864_inst_req_1 : boolean;
  signal type_cast_2194_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1879_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1895_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1910_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1876_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1876_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1882_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1879_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1882_inst_req_0 : boolean;
  signal type_cast_1899_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1861_inst_ack_1 : boolean;
  signal type_cast_1899_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1861_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1858_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1913_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1913_inst_ack_0 : boolean;
  signal type_cast_2029_inst_req_0 : boolean;
  signal type_cast_2029_inst_ack_0 : boolean;
  signal type_cast_1886_inst_ack_1 : boolean;
  signal type_cast_1958_inst_req_1 : boolean;
  signal type_cast_1886_inst_req_1 : boolean;
  signal type_cast_1958_inst_req_0 : boolean;
  signal type_cast_1958_inst_ack_0 : boolean;
  signal type_cast_1958_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1876_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1876_inst_req_0 : boolean;
  signal type_cast_1886_inst_ack_0 : boolean;
  signal type_cast_1954_inst_req_1 : boolean;
  signal type_cast_1954_inst_ack_1 : boolean;
  signal type_cast_1886_inst_req_0 : boolean;
  signal type_cast_1954_inst_req_0 : boolean;
  signal type_cast_1954_inst_ack_0 : boolean;
  signal phi_stmt_2176_req_1 : boolean;
  signal type_cast_1946_inst_req_0 : boolean;
  signal type_cast_1950_inst_req_0 : boolean;
  signal type_cast_1950_inst_ack_0 : boolean;
  signal type_cast_1950_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1861_inst_ack_0 : boolean;
  signal type_cast_1950_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1873_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1882_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1873_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1882_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1861_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1855_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1867_inst_ack_1 : boolean;
  signal type_cast_1946_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1855_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1867_inst_req_1 : boolean;
  signal type_cast_1946_inst_req_1 : boolean;
  signal type_cast_2029_inst_req_1 : boolean;
  signal type_cast_2029_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1855_inst_ack_0 : boolean;
  signal type_cast_2194_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1855_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1907_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1873_inst_ack_0 : boolean;
  signal type_cast_1946_inst_ack_0 : boolean;
  signal type_cast_2033_inst_req_0 : boolean;
  signal type_cast_2033_inst_ack_0 : boolean;
  signal type_cast_2194_inst_ack_1 : boolean;
  signal type_cast_2033_inst_req_1 : boolean;
  signal type_cast_2033_inst_ack_1 : boolean;
  signal type_cast_2037_inst_req_0 : boolean;
  signal type_cast_2037_inst_ack_0 : boolean;
  signal type_cast_2188_inst_req_1 : boolean;
  signal type_cast_2037_inst_req_1 : boolean;
  signal type_cast_2037_inst_ack_1 : boolean;
  signal phi_stmt_2189_ack_0 : boolean;
  signal type_cast_2067_inst_req_0 : boolean;
  signal type_cast_2067_inst_ack_0 : boolean;
  signal type_cast_2067_inst_req_1 : boolean;
  signal type_cast_2067_inst_ack_1 : boolean;
  signal phi_stmt_2183_ack_0 : boolean;
  signal phi_stmt_2176_ack_0 : boolean;
  signal phi_stmt_2189_req_0 : boolean;
  signal type_cast_2192_inst_ack_1 : boolean;
  signal array_obj_ref_2073_index_offset_req_0 : boolean;
  signal array_obj_ref_2073_index_offset_ack_0 : boolean;
  signal array_obj_ref_2073_index_offset_req_1 : boolean;
  signal array_obj_ref_2073_index_offset_ack_1 : boolean;
  signal type_cast_2192_inst_req_1 : boolean;
  signal addr_of_2074_final_reg_req_0 : boolean;
  signal addr_of_2074_final_reg_ack_0 : boolean;
  signal addr_of_2074_final_reg_req_1 : boolean;
  signal addr_of_2074_final_reg_ack_1 : boolean;
  signal type_cast_2192_inst_ack_0 : boolean;
  signal ptr_deref_2078_load_0_req_0 : boolean;
  signal type_cast_2192_inst_req_0 : boolean;
  signal ptr_deref_2078_load_0_ack_0 : boolean;
  signal type_cast_2188_inst_ack_0 : boolean;
  signal ptr_deref_2078_load_0_req_1 : boolean;
  signal ptr_deref_2078_load_0_ack_1 : boolean;
  signal array_obj_ref_2096_index_offset_req_0 : boolean;
  signal array_obj_ref_2096_index_offset_ack_0 : boolean;
  signal array_obj_ref_2096_index_offset_req_1 : boolean;
  signal array_obj_ref_2096_index_offset_ack_1 : boolean;
  signal addr_of_2097_final_reg_req_0 : boolean;
  signal addr_of_2097_final_reg_ack_0 : boolean;
  signal addr_of_2097_final_reg_req_1 : boolean;
  signal addr_of_2097_final_reg_ack_1 : boolean;
  signal phi_stmt_2176_req_0 : boolean;
  signal type_cast_2188_inst_req_0 : boolean;
  signal ptr_deref_2100_store_0_req_0 : boolean;
  signal type_cast_2179_inst_ack_1 : boolean;
  signal ptr_deref_2100_store_0_ack_0 : boolean;
  signal ptr_deref_2100_store_0_req_1 : boolean;
  signal type_cast_2179_inst_req_1 : boolean;
  signal ptr_deref_2100_store_0_ack_1 : boolean;
  signal type_cast_2105_inst_req_0 : boolean;
  signal type_cast_2105_inst_ack_0 : boolean;
  signal type_cast_2105_inst_req_1 : boolean;
  signal type_cast_2105_inst_ack_1 : boolean;
  signal phi_stmt_2183_req_0 : boolean;
  signal if_stmt_2118_branch_req_0 : boolean;
  signal type_cast_2186_inst_ack_1 : boolean;
  signal type_cast_2186_inst_req_1 : boolean;
  signal if_stmt_2118_branch_ack_1 : boolean;
  signal if_stmt_2118_branch_ack_0 : boolean;
  signal type_cast_2186_inst_ack_0 : boolean;
  signal type_cast_2146_inst_req_0 : boolean;
  signal type_cast_2146_inst_ack_0 : boolean;
  signal type_cast_2146_inst_req_1 : boolean;
  signal type_cast_2146_inst_ack_1 : boolean;
  signal type_cast_2179_inst_ack_0 : boolean;
  signal type_cast_2162_inst_req_0 : boolean;
  signal type_cast_2162_inst_ack_0 : boolean;
  signal type_cast_2162_inst_req_1 : boolean;
  signal type_cast_2162_inst_ack_1 : boolean;
  signal type_cast_2179_inst_req_0 : boolean;
  signal type_cast_2186_inst_req_0 : boolean;
  signal if_stmt_2169_branch_req_0 : boolean;
  signal if_stmt_2169_branch_ack_1 : boolean;
  signal if_stmt_2169_branch_ack_0 : boolean;
  signal WPIPE_Block1_done_2205_inst_req_0 : boolean;
  signal WPIPE_Block1_done_2205_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2205_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2205_inst_ack_1 : boolean;
  signal type_cast_1992_inst_req_0 : boolean;
  signal type_cast_1992_inst_ack_0 : boolean;
  signal type_cast_1992_inst_req_1 : boolean;
  signal type_cast_1992_inst_ack_1 : boolean;
  signal phi_stmt_1989_req_0 : boolean;
  signal phi_stmt_1982_req_1 : boolean;
  signal phi_stmt_1975_req_0 : boolean;
  signal phi_stmt_1968_req_0 : boolean;
  signal type_cast_1994_inst_req_0 : boolean;
  signal type_cast_1994_inst_ack_0 : boolean;
  signal type_cast_1994_inst_req_1 : boolean;
  signal type_cast_1994_inst_ack_1 : boolean;
  signal phi_stmt_1989_req_1 : boolean;
  signal type_cast_1985_inst_req_0 : boolean;
  signal type_cast_1985_inst_ack_0 : boolean;
  signal type_cast_1985_inst_req_1 : boolean;
  signal type_cast_1985_inst_ack_1 : boolean;
  signal phi_stmt_1982_req_0 : boolean;
  signal type_cast_1981_inst_req_0 : boolean;
  signal type_cast_1981_inst_ack_0 : boolean;
  signal type_cast_1981_inst_req_1 : boolean;
  signal type_cast_1981_inst_ack_1 : boolean;
  signal phi_stmt_1975_req_1 : boolean;
  signal type_cast_1974_inst_req_0 : boolean;
  signal type_cast_1974_inst_ack_0 : boolean;
  signal type_cast_1974_inst_req_1 : boolean;
  signal phi_stmt_2183_req_1 : boolean;
  signal type_cast_1974_inst_ack_1 : boolean;
  signal phi_stmt_1968_req_1 : boolean;
  signal type_cast_2188_inst_ack_1 : boolean;
  signal phi_stmt_1968_ack_0 : boolean;
  signal phi_stmt_1975_ack_0 : boolean;
  signal phi_stmt_1982_ack_0 : boolean;
  signal phi_stmt_1989_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_4753_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4753_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_4753_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4753_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_4753: Block -- control-path 
    signal convTransposeB_CP_4753_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_4753_elements(0) <= convTransposeB_CP_4753_start;
    convTransposeB_CP_4753_symbol <= convTransposeB_CP_4753_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914__entry__
      -- CP-element group 0: 	 branch_block_stmt_1853/$entry
      -- CP-element group 0: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1855_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1853/branch_block_stmt_1853__entry__
      -- CP-element group 0: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1855_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1899_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1886_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1899_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1899_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1886_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1886_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1855_Sample/rr
      -- 
    cr_4974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(0), ack => type_cast_1899_inst_req_1); -- 
    cr_4946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(0), ack => type_cast_1886_inst_req_1); -- 
    rr_4801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(0), ack => RPIPE_Block1_start_1855_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1853/assign_stmt_2201__exit__
      -- CP-element group 1: 	 branch_block_stmt_1853/assign_stmt_2201__entry__
      -- CP-element group 1: 	 branch_block_stmt_1853/merge_stmt_2175__exit__
      -- CP-element group 1: 	 branch_block_stmt_1853/assign_stmt_2201/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/assign_stmt_2201/$exit
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1989/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1994/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1994/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1994/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1994/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1994/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1994/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1982/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_sources/type_cast_1985/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_sources/type_cast_1985/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_sources/type_cast_1985/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_sources/type_cast_1985/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_sources/type_cast_1985/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_sources/type_cast_1985/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1975/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_sources/type_cast_1981/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_sources/type_cast_1981/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_sources/type_cast_1981/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_sources/type_cast_1981/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_sources/type_cast_1981/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_sources/type_cast_1981/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1968/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_sources/type_cast_1974/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_sources/type_cast_1974/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_sources/type_cast_1974/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_sources/type_cast_1974/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_sources/type_cast_1974/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_sources/type_cast_1974/SplitProtocol/Update/cr
      -- 
    rr_5502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(1), ack => type_cast_1994_inst_req_0); -- 
    cr_5507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(1), ack => type_cast_1994_inst_req_1); -- 
    rr_5525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(1), ack => type_cast_1985_inst_req_0); -- 
    cr_5530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(1), ack => type_cast_1985_inst_req_1); -- 
    rr_5548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(1), ack => type_cast_1981_inst_req_0); -- 
    cr_5553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(1), ack => type_cast_1981_inst_req_1); -- 
    rr_5571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(1), ack => type_cast_1974_inst_req_0); -- 
    cr_5576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(1), ack => type_cast_1974_inst_req_1); -- 
    convTransposeB_CP_4753_elements(1) <= convTransposeB_CP_4753_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1855_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1855_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1855_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1855_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1855_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1855_Sample/$exit
      -- 
    ra_4802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1855_inst_ack_0, ack => convTransposeB_CP_4753_elements(2)); -- 
    cr_4806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(2), ack => RPIPE_Block1_start_1855_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1858_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1855_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1858_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1858_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1855_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1855_Update/$exit
      -- 
    ca_4807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1855_inst_ack_1, ack => convTransposeB_CP_4753_elements(3)); -- 
    rr_4815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(3), ack => RPIPE_Block1_start_1858_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1858_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1858_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1858_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1858_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1858_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1858_sample_completed_
      -- 
    ra_4816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1858_inst_ack_0, ack => convTransposeB_CP_4753_elements(4)); -- 
    cr_4820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(4), ack => RPIPE_Block1_start_1858_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1858_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1858_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1858_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1861_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1861_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1861_Sample/$entry
      -- 
    ca_4821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1858_inst_ack_1, ack => convTransposeB_CP_4753_elements(5)); -- 
    rr_4829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(5), ack => RPIPE_Block1_start_1861_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1861_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1861_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1861_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1861_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1861_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1861_Sample/$exit
      -- 
    ra_4830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1861_inst_ack_0, ack => convTransposeB_CP_4753_elements(6)); -- 
    cr_4834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(6), ack => RPIPE_Block1_start_1861_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1864_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1864_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1864_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1861_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1861_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1861_update_completed_
      -- 
    ca_4835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1861_inst_ack_1, ack => convTransposeB_CP_4753_elements(7)); -- 
    rr_4843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(7), ack => RPIPE_Block1_start_1864_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1864_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1864_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1864_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1864_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1864_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1864_sample_completed_
      -- 
    ra_4844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1864_inst_ack_0, ack => convTransposeB_CP_4753_elements(8)); -- 
    cr_4848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(8), ack => RPIPE_Block1_start_1864_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1867_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1864_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1864_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1867_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1867_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1864_Update/$exit
      -- 
    ca_4849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1864_inst_ack_1, ack => convTransposeB_CP_4753_elements(9)); -- 
    rr_4857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(9), ack => RPIPE_Block1_start_1867_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1867_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1867_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1867_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1867_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1867_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1867_Update/cr
      -- 
    ra_4858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1867_inst_ack_0, ack => convTransposeB_CP_4753_elements(10)); -- 
    cr_4862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(10), ack => RPIPE_Block1_start_1867_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1870_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1870_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1867_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1870_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1867_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1867_Update/$exit
      -- 
    ca_4863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1867_inst_ack_1, ack => convTransposeB_CP_4753_elements(11)); -- 
    rr_4871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(11), ack => RPIPE_Block1_start_1870_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1870_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1870_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1870_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1870_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1870_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1870_sample_completed_
      -- 
    ra_4872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1870_inst_ack_0, ack => convTransposeB_CP_4753_elements(12)); -- 
    cr_4876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(12), ack => RPIPE_Block1_start_1870_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1870_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1873_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1870_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1873_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1873_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1870_update_completed_
      -- 
    ca_4877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1870_inst_ack_1, ack => convTransposeB_CP_4753_elements(13)); -- 
    rr_4885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(13), ack => RPIPE_Block1_start_1873_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1873_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1873_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1873_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1873_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1873_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1873_Sample/ra
      -- 
    ra_4886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1873_inst_ack_0, ack => convTransposeB_CP_4753_elements(14)); -- 
    cr_4890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(14), ack => RPIPE_Block1_start_1873_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1873_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1876_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1876_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1876_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1873_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1873_Update/$exit
      -- 
    ca_4891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1873_inst_ack_1, ack => convTransposeB_CP_4753_elements(15)); -- 
    rr_4899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(15), ack => RPIPE_Block1_start_1876_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1876_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1876_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1876_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1876_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1876_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1876_sample_completed_
      -- 
    ra_4900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1876_inst_ack_0, ack => convTransposeB_CP_4753_elements(16)); -- 
    cr_4904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(16), ack => RPIPE_Block1_start_1876_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1879_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1879_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1879_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1876_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1876_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1876_update_completed_
      -- 
    ca_4905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1876_inst_ack_1, ack => convTransposeB_CP_4753_elements(17)); -- 
    rr_4913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(17), ack => RPIPE_Block1_start_1879_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1879_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1879_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1879_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1879_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1879_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1879_Update/cr
      -- 
    ra_4914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1879_inst_ack_0, ack => convTransposeB_CP_4753_elements(18)); -- 
    cr_4918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(18), ack => RPIPE_Block1_start_1879_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1879_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1879_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1879_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1882_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1882_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1882_sample_start_
      -- 
    ca_4919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1879_inst_ack_1, ack => convTransposeB_CP_4753_elements(19)); -- 
    rr_4927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(19), ack => RPIPE_Block1_start_1882_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1882_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1882_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1882_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1882_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1882_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1882_sample_completed_
      -- 
    ra_4928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1882_inst_ack_0, ack => convTransposeB_CP_4753_elements(20)); -- 
    cr_4932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(20), ack => RPIPE_Block1_start_1882_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1882_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1895_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1895_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1895_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1886_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1886_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1886_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1882_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1882_update_completed_
      -- 
    ca_4933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1882_inst_ack_1, ack => convTransposeB_CP_4753_elements(21)); -- 
    rr_4941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(21), ack => type_cast_1886_inst_req_0); -- 
    rr_4955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(21), ack => RPIPE_Block1_start_1895_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1886_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1886_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1886_sample_completed_
      -- 
    ra_4942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1886_inst_ack_0, ack => convTransposeB_CP_4753_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1886_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1886_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1886_update_completed_
      -- 
    ca_4947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1886_inst_ack_1, ack => convTransposeB_CP_4753_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1895_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1895_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1895_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1895_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1895_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1895_sample_completed_
      -- 
    ra_4956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1895_inst_ack_0, ack => convTransposeB_CP_4753_elements(24)); -- 
    cr_4960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(24), ack => RPIPE_Block1_start_1895_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1895_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1899_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1899_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1895_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1907_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1907_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1895_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1907_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1899_sample_start_
      -- 
    ca_4961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1895_inst_ack_1, ack => convTransposeB_CP_4753_elements(25)); -- 
    rr_4969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(25), ack => type_cast_1899_inst_req_0); -- 
    rr_4983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(25), ack => RPIPE_Block1_start_1907_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1899_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1899_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1899_Sample/ra
      -- 
    ra_4970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1899_inst_ack_0, ack => convTransposeB_CP_4753_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1899_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1899_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/type_cast_1899_Update/$exit
      -- 
    ca_4975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1899_inst_ack_1, ack => convTransposeB_CP_4753_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1907_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1907_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1907_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1907_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1907_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1907_sample_completed_
      -- 
    ra_4984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1907_inst_ack_0, ack => convTransposeB_CP_4753_elements(28)); -- 
    cr_4988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(28), ack => RPIPE_Block1_start_1907_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1910_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1907_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1907_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1910_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1907_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1910_Sample/$entry
      -- 
    ca_4989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1907_inst_ack_1, ack => convTransposeB_CP_4753_elements(29)); -- 
    rr_4997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(29), ack => RPIPE_Block1_start_1910_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1910_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1910_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1910_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1910_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1910_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1910_sample_completed_
      -- 
    ra_4998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1910_inst_ack_0, ack => convTransposeB_CP_4753_elements(30)); -- 
    cr_5002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(30), ack => RPIPE_Block1_start_1910_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1913_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1910_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1913_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1910_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1913_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1910_update_completed_
      -- 
    ca_5003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1910_inst_ack_1, ack => convTransposeB_CP_4753_elements(31)); -- 
    rr_5011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(31), ack => RPIPE_Block1_start_1913_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1913_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1913_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1913_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1913_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1913_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1913_Sample/ra
      -- 
    ra_5012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1913_inst_ack_0, ack => convTransposeB_CP_4753_elements(32)); -- 
    cr_5016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(32), ack => RPIPE_Block1_start_1913_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1913_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1913_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/RPIPE_Block1_start_1913_Update/$exit
      -- 
    ca_5017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1913_inst_ack_1, ack => convTransposeB_CP_4753_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914/$exit
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1856_to_assign_stmt_1914__exit__
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965__entry__
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1958_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1958_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1958_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1958_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1958_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1958_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1954_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1954_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1954_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1954_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1954_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1954_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1946_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1946_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1950_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1950_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1950_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1950_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1950_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1950_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1946_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1946_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/$entry
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1946_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1946_update_start_
      -- 
    cr_5075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(34), ack => type_cast_1958_inst_req_1); -- 
    rr_5070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(34), ack => type_cast_1958_inst_req_0); -- 
    cr_5061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(34), ack => type_cast_1954_inst_req_1); -- 
    rr_5056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(34), ack => type_cast_1954_inst_req_0); -- 
    rr_5028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(34), ack => type_cast_1946_inst_req_0); -- 
    rr_5042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(34), ack => type_cast_1950_inst_req_0); -- 
    cr_5047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(34), ack => type_cast_1950_inst_req_1); -- 
    cr_5033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(34), ack => type_cast_1946_inst_req_1); -- 
    convTransposeB_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(23) & convTransposeB_CP_4753_elements(27) & convTransposeB_CP_4753_elements(33);
      gj_convTransposeB_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1946_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1946_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1946_Sample/ra
      -- 
    ra_5029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1946_inst_ack_0, ack => convTransposeB_CP_4753_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1946_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1946_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1946_update_completed_
      -- 
    ca_5034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1946_inst_ack_1, ack => convTransposeB_CP_4753_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1950_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1950_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1950_sample_completed_
      -- 
    ra_5043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1950_inst_ack_0, ack => convTransposeB_CP_4753_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1950_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1950_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1950_update_completed_
      -- 
    ca_5048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1950_inst_ack_1, ack => convTransposeB_CP_4753_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1954_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1954_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1954_sample_completed_
      -- 
    ra_5057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1954_inst_ack_0, ack => convTransposeB_CP_4753_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1954_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1954_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1954_update_completed_
      -- 
    ca_5062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1954_inst_ack_1, ack => convTransposeB_CP_4753_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1958_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1958_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1958_sample_completed_
      -- 
    ra_5071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1958_inst_ack_0, ack => convTransposeB_CP_4753_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1958_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1958_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/type_cast_1958_update_completed_
      -- 
    ca_5076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1958_inst_ack_1, ack => convTransposeB_CP_4753_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	82 
    -- CP-element group 43: 	83 
    -- CP-element group 43: 	84 
    -- CP-element group 43:  members (18) 
      -- CP-element group 43: 	 branch_block_stmt_1853/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965__exit__
      -- CP-element group 43: 	 branch_block_stmt_1853/assign_stmt_1921_to_assign_stmt_1965/$exit
      -- CP-element group 43: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1989/$entry
      -- CP-element group 43: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1992/$entry
      -- CP-element group 43: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1992/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1992/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1992/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1992/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1992/SplitProtocol/Update/cr
      -- CP-element group 43: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1982/$entry
      -- CP-element group 43: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1975/$entry
      -- CP-element group 43: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1968/$entry
      -- CP-element group 43: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_sources/$entry
      -- 
    rr_5452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(43), ack => type_cast_1992_inst_req_0); -- 
    cr_5457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(43), ack => type_cast_1992_inst_req_1); -- 
    convTransposeB_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(36) & convTransposeB_CP_4753_elements(38) & convTransposeB_CP_4753_elements(40) & convTransposeB_CP_4753_elements(42);
      gj_convTransposeB_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	104 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2029_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2029_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2029_Sample/$exit
      -- 
    ra_5088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2029_inst_ack_0, ack => convTransposeB_CP_4753_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	104 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2029_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2029_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2029_Update/ca
      -- 
    ca_5093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2029_inst_ack_1, ack => convTransposeB_CP_4753_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	104 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2033_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2033_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2033_Sample/ra
      -- 
    ra_5102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2033_inst_ack_0, ack => convTransposeB_CP_4753_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	104 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2033_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2033_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2033_Update/ca
      -- 
    ca_5107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2033_inst_ack_1, ack => convTransposeB_CP_4753_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	104 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2037_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2037_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2037_Sample/ra
      -- 
    ra_5116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2037_inst_ack_0, ack => convTransposeB_CP_4753_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	104 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2037_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2037_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2037_Update/ca
      -- 
    ca_5121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2037_inst_ack_1, ack => convTransposeB_CP_4753_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	104 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2067_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2067_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2067_Sample/ra
      -- 
    ra_5130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2067_inst_ack_0, ack => convTransposeB_CP_4753_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	104 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2067_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2067_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2067_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_final_index_sum_regn_Sample/req
      -- 
    ca_5135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2067_inst_ack_1, ack => convTransposeB_CP_4753_elements(51)); -- 
    req_5160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(51), ack => array_obj_ref_2073_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_final_index_sum_regn_Sample/ack
      -- 
    ack_5161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2073_index_offset_ack_0, ack => convTransposeB_CP_4753_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	104 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2074_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2074_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2074_request/req
      -- 
    ack_5166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2073_index_offset_ack_1, ack => convTransposeB_CP_4753_elements(53)); -- 
    req_5175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(53), ack => addr_of_2074_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2074_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2074_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2074_request/ack
      -- 
    ack_5176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2074_final_reg_ack_0, ack => convTransposeB_CP_4753_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	104 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2074_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2074_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2074_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Sample/word_access_start/word_0/rr
      -- 
    ack_5181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2074_final_reg_ack_1, ack => convTransposeB_CP_4753_elements(55)); -- 
    rr_5214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(55), ack => ptr_deref_2078_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Sample/word_access_start/word_0/ra
      -- 
    ra_5215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2078_load_0_ack_0, ack => convTransposeB_CP_4753_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	104 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Update/ptr_deref_2078_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Update/ptr_deref_2078_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Update/ptr_deref_2078_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Update/ptr_deref_2078_Merge/merge_ack
      -- 
    ca_5226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2078_load_0_ack_1, ack => convTransposeB_CP_4753_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_final_index_sum_regn_Sample/req
      -- 
    req_5256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(58), ack => array_obj_ref_2096_index_offset_req_0); -- 
    convTransposeB_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(45) & convTransposeB_CP_4753_elements(47) & convTransposeB_CP_4753_elements(49);
      gj_convTransposeB_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_final_index_sum_regn_Sample/ack
      -- 
    ack_5257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2096_index_offset_ack_0, ack => convTransposeB_CP_4753_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	104 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2097_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2097_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2097_request/req
      -- 
    ack_5262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2096_index_offset_ack_1, ack => convTransposeB_CP_4753_elements(60)); -- 
    req_5271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(60), ack => addr_of_2097_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2097_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2097_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2097_request/ack
      -- 
    ack_5272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2097_final_reg_ack_0, ack => convTransposeB_CP_4753_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	104 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2097_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2097_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2097_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_word_addrgen/root_register_ack
      -- 
    ack_5277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2097_final_reg_ack_1, ack => convTransposeB_CP_4753_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Sample/ptr_deref_2100_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Sample/ptr_deref_2100_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Sample/ptr_deref_2100_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Sample/ptr_deref_2100_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Sample/word_access_start/word_0/rr
      -- 
    rr_5315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(63), ack => ptr_deref_2100_store_0_req_0); -- 
    convTransposeB_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(57) & convTransposeB_CP_4753_elements(62);
      gj_convTransposeB_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Sample/word_access_start/word_0/ra
      -- 
    ra_5316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2100_store_0_ack_0, ack => convTransposeB_CP_4753_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	104 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Update/word_access_complete/word_0/ca
      -- 
    ca_5327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2100_store_0_ack_1, ack => convTransposeB_CP_4753_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	104 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2105_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2105_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2105_Sample/ra
      -- 
    ra_5336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2105_inst_ack_0, ack => convTransposeB_CP_4753_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	104 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2105_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2105_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2105_Update/ca
      -- 
    ca_5341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2105_inst_ack_1, ack => convTransposeB_CP_4753_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117__exit__
      -- CP-element group 68: 	 branch_block_stmt_1853/if_stmt_2118__entry__
      -- CP-element group 68: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/$exit
      -- CP-element group 68: 	 branch_block_stmt_1853/if_stmt_2118_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1853/if_stmt_2118_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1853/if_stmt_2118_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1853/if_stmt_2118_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1853/R_cmp_2119_place
      -- CP-element group 68: 	 branch_block_stmt_1853/if_stmt_2118_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1853/if_stmt_2118_else_link/$entry
      -- 
    branch_req_5349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(68), ack => if_stmt_2118_branch_req_0); -- 
    convTransposeB_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(52) & convTransposeB_CP_4753_elements(59) & convTransposeB_CP_4753_elements(65) & convTransposeB_CP_4753_elements(67);
      gj_convTransposeB_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	113 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	116 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	119 
    -- CP-element group 69: 	120 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_1853/assign_stmt_2130__entry__
      -- CP-element group 69: 	 branch_block_stmt_1853/merge_stmt_2124__exit__
      -- CP-element group 69: 	 branch_block_stmt_1853/assign_stmt_2130__exit__
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2192/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2192/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2192/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2192/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2192/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2192/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2189/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_sources/type_cast_2179/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_sources/type_cast_2179/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/if_stmt_2118_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1853/if_stmt_2118_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1853/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_1853/assign_stmt_2130/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/assign_stmt_2130/$exit
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_sources/type_cast_2179/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_sources/type_cast_2179/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_sources/type_cast_2179/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_sources/type_cast_2179/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2176/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1853/merge_stmt_2124_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1853/merge_stmt_2124_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1853/merge_stmt_2124_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1853/merge_stmt_2124_PhiAck/dummy
      -- 
    if_choice_transition_5354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2118_branch_ack_1, ack => convTransposeB_CP_4753_elements(69)); -- 
    cr_5691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(69), ack => type_cast_2188_inst_req_1); -- 
    cr_5737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(69), ack => type_cast_2192_inst_req_1); -- 
    rr_5732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(69), ack => type_cast_2192_inst_req_0); -- 
    rr_5686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(69), ack => type_cast_2188_inst_req_0); -- 
    cr_5714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(69), ack => type_cast_2179_inst_req_1); -- 
    rr_5709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(69), ack => type_cast_2179_inst_req_0); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_1853/merge_stmt_2132__exit__
      -- CP-element group 70: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168__entry__
      -- CP-element group 70: 	 branch_block_stmt_1853/if_stmt_2118_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1853/if_stmt_2118_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1853/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/$entry
      -- CP-element group 70: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2146_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2146_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2146_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2146_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2146_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2146_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2162_update_start_
      -- CP-element group 70: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2162_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2162_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1853/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1853/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_1853/merge_stmt_2132_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_1853/merge_stmt_2132_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_1853/merge_stmt_2132_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_1853/merge_stmt_2132_PhiAck/dummy
      -- 
    else_choice_transition_5358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2118_branch_ack_0, ack => convTransposeB_CP_4753_elements(70)); -- 
    rr_5374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(70), ack => type_cast_2146_inst_req_0); -- 
    cr_5379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(70), ack => type_cast_2146_inst_req_1); -- 
    cr_5393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(70), ack => type_cast_2162_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2146_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2146_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2146_Sample/ra
      -- 
    ra_5375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2146_inst_ack_0, ack => convTransposeB_CP_4753_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2146_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2146_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2146_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2162_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2162_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2162_Sample/rr
      -- 
    ca_5380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2146_inst_ack_1, ack => convTransposeB_CP_4753_elements(72)); -- 
    rr_5388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(72), ack => type_cast_2162_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2162_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2162_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2162_Sample/ra
      -- 
    ra_5389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2162_inst_ack_0, ack => convTransposeB_CP_4753_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_1853/if_stmt_2169__entry__
      -- CP-element group 74: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168__exit__
      -- CP-element group 74: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/$exit
      -- CP-element group 74: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2162_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2162_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1853/assign_stmt_2138_to_assign_stmt_2168/type_cast_2162_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_1853/if_stmt_2169_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1853/if_stmt_2169_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_1853/if_stmt_2169_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_1853/if_stmt_2169_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_1853/R_cmp117_2170_place
      -- CP-element group 74: 	 branch_block_stmt_1853/if_stmt_2169_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_1853/if_stmt_2169_else_link/$entry
      -- 
    ca_5394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2162_inst_ack_1, ack => convTransposeB_CP_4753_elements(74)); -- 
    branch_req_5402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(74), ack => if_stmt_2169_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_1853/merge_stmt_2203__exit__
      -- CP-element group 75: 	 branch_block_stmt_1853/assign_stmt_2208__entry__
      -- CP-element group 75: 	 branch_block_stmt_1853/merge_stmt_2203_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_1853/merge_stmt_2203_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_1853/merge_stmt_2203_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_1853/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_1853/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_1853/merge_stmt_2203_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_1853/if_stmt_2169_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_1853/if_stmt_2169_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_1853/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_1853/assign_stmt_2208/$entry
      -- CP-element group 75: 	 branch_block_stmt_1853/assign_stmt_2208/WPIPE_Block1_done_2205_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1853/assign_stmt_2208/WPIPE_Block1_done_2205_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1853/assign_stmt_2208/WPIPE_Block1_done_2205_Sample/req
      -- 
    if_choice_transition_5407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2169_branch_ack_1, ack => convTransposeB_CP_4753_elements(75)); -- 
    req_5427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(75), ack => WPIPE_Block1_done_2205_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	108 
    -- CP-element group 76: 	109 
    -- CP-element group 76: 	110 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2194/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2194/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/$entry
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2194/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2189/$entry
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2194/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2194/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2176/$entry
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_1853/if_stmt_2169_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_1853/if_stmt_2169_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/$entry
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2194/$entry
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/$entry
      -- 
    else_choice_transition_5411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2169_branch_ack_0, ack => convTransposeB_CP_4753_elements(76)); -- 
    rr_5660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(76), ack => type_cast_2194_inst_req_0); -- 
    cr_5665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(76), ack => type_cast_2194_inst_req_1); -- 
    cr_5634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(76), ack => type_cast_2186_inst_req_1); -- 
    rr_5629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(76), ack => type_cast_2186_inst_req_0); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_1853/assign_stmt_2208/WPIPE_Block1_done_2205_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1853/assign_stmt_2208/WPIPE_Block1_done_2205_update_start_
      -- CP-element group 77: 	 branch_block_stmt_1853/assign_stmt_2208/WPIPE_Block1_done_2205_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1853/assign_stmt_2208/WPIPE_Block1_done_2205_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_1853/assign_stmt_2208/WPIPE_Block1_done_2205_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_1853/assign_stmt_2208/WPIPE_Block1_done_2205_Update/req
      -- 
    ack_5428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2205_inst_ack_0, ack => convTransposeB_CP_4753_elements(77)); -- 
    req_5432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(77), ack => WPIPE_Block1_done_2205_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 branch_block_stmt_1853/branch_block_stmt_1853__exit__
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_1853/assign_stmt_2208__exit__
      -- CP-element group 78: 	 branch_block_stmt_1853/return__
      -- CP-element group 78: 	 branch_block_stmt_1853/$exit
      -- CP-element group 78: 	 branch_block_stmt_1853/merge_stmt_2210__exit__
      -- CP-element group 78: 	 branch_block_stmt_1853/merge_stmt_2210_PhiAck/dummy
      -- CP-element group 78: 	 branch_block_stmt_1853/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_1853/merge_stmt_2210_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_1853/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_1853/merge_stmt_2210_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_1853/merge_stmt_2210_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_1853/assign_stmt_2208/$exit
      -- CP-element group 78: 	 branch_block_stmt_1853/assign_stmt_2208/WPIPE_Block1_done_2205_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1853/assign_stmt_2208/WPIPE_Block1_done_2205_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1853/assign_stmt_2208/WPIPE_Block1_done_2205_Update/ack
      -- 
    ack_5433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2205_inst_ack_1, ack => convTransposeB_CP_4753_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1992/SplitProtocol/Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1992/SplitProtocol/Sample/ra
      -- 
    ra_5453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1992_inst_ack_0, ack => convTransposeB_CP_4753_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1992/SplitProtocol/Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1992/SplitProtocol/Update/ca
      -- 
    ca_5458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1992_inst_ack_1, ack => convTransposeB_CP_4753_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1989/$exit
      -- CP-element group 81: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1992/$exit
      -- CP-element group 81: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1992/SplitProtocol/$exit
      -- CP-element group 81: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_req
      -- 
    phi_stmt_1989_req_5459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1989_req_5459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(81), ack => phi_stmt_1989_req_0); -- 
    convTransposeB_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(79) & convTransposeB_CP_4753_elements(80);
      gj_convTransposeB_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  output  delay-element  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	85 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1982/$exit
      -- CP-element group 82: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_sources/type_cast_1988_konst_delay_trans
      -- CP-element group 82: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_req
      -- 
    phi_stmt_1982_req_5467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1982_req_5467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(82), ack => phi_stmt_1982_req_1); -- 
    -- Element group convTransposeB_CP_4753_elements(82) is a control-delay.
    cp_element_82_delay: control_delay_element  generic map(name => " 82_delay", delay_value => 1)  port map(req => convTransposeB_CP_4753_elements(43), ack => convTransposeB_CP_4753_elements(82), clk => clk, reset =>reset);
    -- CP-element group 83:  transition  output  delay-element  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	43 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1975/$exit
      -- CP-element group 83: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_sources/$exit
      -- CP-element group 83: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_sources/type_cast_1979_konst_delay_trans
      -- CP-element group 83: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_req
      -- 
    phi_stmt_1975_req_5475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1975_req_5475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(83), ack => phi_stmt_1975_req_0); -- 
    -- Element group convTransposeB_CP_4753_elements(83) is a control-delay.
    cp_element_83_delay: control_delay_element  generic map(name => " 83_delay", delay_value => 1)  port map(req => convTransposeB_CP_4753_elements(43), ack => convTransposeB_CP_4753_elements(83), clk => clk, reset =>reset);
    -- CP-element group 84:  transition  output  delay-element  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	43 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1968/$exit
      -- CP-element group 84: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_sources/type_cast_1972_konst_delay_trans
      -- CP-element group 84: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_req
      -- 
    phi_stmt_1968_req_5483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1968_req_5483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(84), ack => phi_stmt_1968_req_0); -- 
    -- Element group convTransposeB_CP_4753_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => convTransposeB_CP_4753_elements(43), ack => convTransposeB_CP_4753_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	81 
    -- CP-element group 85: 	82 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	99 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1853/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(81) & convTransposeB_CP_4753_elements(82) & convTransposeB_CP_4753_elements(83) & convTransposeB_CP_4753_elements(84);
      gj_convTransposeB_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1994/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1994/SplitProtocol/Sample/ra
      -- 
    ra_5503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1994_inst_ack_0, ack => convTransposeB_CP_4753_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1994/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1994/SplitProtocol/Update/ca
      -- 
    ca_5508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1994_inst_ack_1, ack => convTransposeB_CP_4753_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	98 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1989/$exit
      -- CP-element group 88: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1994/$exit
      -- CP-element group 88: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_sources/type_cast_1994/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1989/phi_stmt_1989_req
      -- 
    phi_stmt_1989_req_5509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1989_req_5509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(88), ack => phi_stmt_1989_req_1); -- 
    convTransposeB_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(86) & convTransposeB_CP_4753_elements(87);
      gj_convTransposeB_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_sources/type_cast_1985/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_sources/type_cast_1985/SplitProtocol/Sample/ra
      -- 
    ra_5526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1985_inst_ack_0, ack => convTransposeB_CP_4753_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_sources/type_cast_1985/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_sources/type_cast_1985/SplitProtocol/Update/ca
      -- 
    ca_5531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1985_inst_ack_1, ack => convTransposeB_CP_4753_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1982/$exit
      -- CP-element group 91: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_sources/type_cast_1985/$exit
      -- CP-element group 91: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_sources/type_cast_1985/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1982/phi_stmt_1982_req
      -- 
    phi_stmt_1982_req_5532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1982_req_5532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(91), ack => phi_stmt_1982_req_0); -- 
    convTransposeB_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(89) & convTransposeB_CP_4753_elements(90);
      gj_convTransposeB_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_sources/type_cast_1981/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_sources/type_cast_1981/SplitProtocol/Sample/ra
      -- 
    ra_5549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1981_inst_ack_0, ack => convTransposeB_CP_4753_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_sources/type_cast_1981/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_sources/type_cast_1981/SplitProtocol/Update/ca
      -- 
    ca_5554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1981_inst_ack_1, ack => convTransposeB_CP_4753_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1975/$exit
      -- CP-element group 94: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_sources/type_cast_1981/$exit
      -- CP-element group 94: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_sources/type_cast_1981/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1975/phi_stmt_1975_req
      -- 
    phi_stmt_1975_req_5555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1975_req_5555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(94), ack => phi_stmt_1975_req_1); -- 
    convTransposeB_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(92) & convTransposeB_CP_4753_elements(93);
      gj_convTransposeB_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_sources/type_cast_1974/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_sources/type_cast_1974/SplitProtocol/Sample/ra
      -- 
    ra_5572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1974_inst_ack_0, ack => convTransposeB_CP_4753_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_sources/type_cast_1974/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_sources/type_cast_1974/SplitProtocol/Update/ca
      -- 
    ca_5577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1974_inst_ack_1, ack => convTransposeB_CP_4753_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1968/$exit
      -- CP-element group 97: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_sources/type_cast_1974/$exit
      -- CP-element group 97: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_sources/type_cast_1974/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/phi_stmt_1968/phi_stmt_1968_req
      -- 
    phi_stmt_1968_req_5578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1968_req_5578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(97), ack => phi_stmt_1968_req_1); -- 
    convTransposeB_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(95) & convTransposeB_CP_4753_elements(96);
      gj_convTransposeB_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1853/ifx_xend128_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(88) & convTransposeB_CP_4753_elements(91) & convTransposeB_CP_4753_elements(94) & convTransposeB_CP_4753_elements(97);
      gj_convTransposeB_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  fork  transition  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	85 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	102 
    -- CP-element group 99: 	103 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1853/merge_stmt_1967_PhiReqMerge
      -- CP-element group 99: 	 branch_block_stmt_1853/merge_stmt_1967_PhiAck/$entry
      -- 
    convTransposeB_CP_4753_elements(99) <= OrReduce(convTransposeB_CP_4753_elements(85) & convTransposeB_CP_4753_elements(98));
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1853/merge_stmt_1967_PhiAck/phi_stmt_1968_ack
      -- 
    phi_stmt_1968_ack_5583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1968_ack_0, ack => convTransposeB_CP_4753_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1853/merge_stmt_1967_PhiAck/phi_stmt_1975_ack
      -- 
    phi_stmt_1975_ack_5584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1975_ack_0, ack => convTransposeB_CP_4753_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1853/merge_stmt_1967_PhiAck/phi_stmt_1982_ack
      -- 
    phi_stmt_1982_ack_5585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1982_ack_0, ack => convTransposeB_CP_4753_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1853/merge_stmt_1967_PhiAck/phi_stmt_1989_ack
      -- 
    phi_stmt_1989_ack_5586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1989_ack_0, ack => convTransposeB_CP_4753_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	44 
    -- CP-element group 104: 	45 
    -- CP-element group 104: 	46 
    -- CP-element group 104: 	47 
    -- CP-element group 104: 	48 
    -- CP-element group 104: 	49 
    -- CP-element group 104: 	50 
    -- CP-element group 104: 	51 
    -- CP-element group 104: 	53 
    -- CP-element group 104: 	55 
    -- CP-element group 104: 	57 
    -- CP-element group 104: 	60 
    -- CP-element group 104: 	62 
    -- CP-element group 104: 	65 
    -- CP-element group 104: 	66 
    -- CP-element group 104: 	67 
    -- CP-element group 104:  members (56) 
      -- CP-element group 104: 	 branch_block_stmt_1853/merge_stmt_1967__exit__
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117__entry__
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2029_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2029_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2029_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2029_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2029_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2029_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2033_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2033_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2033_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2033_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2033_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2033_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2037_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2037_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2037_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2037_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2037_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2037_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2067_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2067_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2067_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2067_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2067_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2067_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2074_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2073_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2074_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2074_complete/req
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2078_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2097_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/array_obj_ref_2096_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2097_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/addr_of_2097_complete/req
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/ptr_deref_2100_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2105_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2105_update_start_
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2105_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2105_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2105_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_1853/assign_stmt_2001_to_assign_stmt_2117/type_cast_2105_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_1853/merge_stmt_1967_PhiAck/$exit
      -- 
    rr_5087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2029_inst_req_0); -- 
    cr_5092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2029_inst_req_1); -- 
    rr_5101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2033_inst_req_0); -- 
    cr_5106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2033_inst_req_1); -- 
    rr_5115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2037_inst_req_0); -- 
    cr_5120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2037_inst_req_1); -- 
    rr_5129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2067_inst_req_0); -- 
    cr_5134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2067_inst_req_1); -- 
    req_5165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => array_obj_ref_2073_index_offset_req_1); -- 
    req_5180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => addr_of_2074_final_reg_req_1); -- 
    cr_5225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => ptr_deref_2078_load_0_req_1); -- 
    req_5261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => array_obj_ref_2096_index_offset_req_1); -- 
    req_5276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => addr_of_2097_final_reg_req_1); -- 
    cr_5326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => ptr_deref_2100_store_0_req_1); -- 
    rr_5335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2105_inst_req_0); -- 
    cr_5340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(104), ack => type_cast_2105_inst_req_1); -- 
    convTransposeB_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(100) & convTransposeB_CP_4753_elements(101) & convTransposeB_CP_4753_elements(102) & convTransposeB_CP_4753_elements(103);
      gj_convTransposeB_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/Sample/$exit
      -- 
    ra_5630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2186_inst_ack_0, ack => convTransposeB_CP_4753_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/Update/ca
      -- CP-element group 106: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/Update/$exit
      -- 
    ca_5635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2186_inst_ack_1, ack => convTransposeB_CP_4753_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	112 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_req
      -- CP-element group 107: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/$exit
      -- CP-element group 107: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2186/$exit
      -- 
    phi_stmt_2183_req_5636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2183_req_5636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(107), ack => phi_stmt_2183_req_0); -- 
    convTransposeB_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(105) & convTransposeB_CP_4753_elements(106);
      gj_convTransposeB_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  transition  output  delay-element  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	76 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_req
      -- CP-element group 108: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_sources/type_cast_2182_konst_delay_trans
      -- CP-element group 108: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2176/$exit
      -- 
    phi_stmt_2176_req_5644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2176_req_5644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(108), ack => phi_stmt_2176_req_1); -- 
    -- Element group convTransposeB_CP_4753_elements(108) is a control-delay.
    cp_element_108_delay: control_delay_element  generic map(name => " 108_delay", delay_value => 1)  port map(req => convTransposeB_CP_4753_elements(76), ack => convTransposeB_CP_4753_elements(108), clk => clk, reset =>reset);
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2194/SplitProtocol/Sample/ra
      -- CP-element group 109: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2194/SplitProtocol/Sample/$exit
      -- 
    ra_5661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2194_inst_ack_0, ack => convTransposeB_CP_4753_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	76 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2194/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2194/SplitProtocol/Update/ca
      -- 
    ca_5666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2194_inst_ack_1, ack => convTransposeB_CP_4753_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_req
      -- CP-element group 111: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2189/$exit
      -- CP-element group 111: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2194/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2194/$exit
      -- CP-element group 111: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/$exit
      -- 
    phi_stmt_2189_req_5667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2189_req_5667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(111), ack => phi_stmt_2189_req_1); -- 
    convTransposeB_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(109) & convTransposeB_CP_4753_elements(110);
      gj_convTransposeB_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	107 
    -- CP-element group 112: 	108 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	123 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1853/ifx_xelse_ifx_xend128_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(107) & convTransposeB_CP_4753_elements(108) & convTransposeB_CP_4753_elements(111);
      gj_convTransposeB_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	69 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/Sample/ra
      -- CP-element group 113: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/Sample/$exit
      -- 
    ra_5687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2188_inst_ack_0, ack => convTransposeB_CP_4753_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/Update/ca
      -- 
    ca_5692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2188_inst_ack_1, ack => convTransposeB_CP_4753_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/type_cast_2188/$exit
      -- CP-element group 115: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/$exit
      -- CP-element group 115: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2183/phi_stmt_2183_req
      -- 
    phi_stmt_2183_req_5693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2183_req_5693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(115), ack => phi_stmt_2183_req_1); -- 
    convTransposeB_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(113) & convTransposeB_CP_4753_elements(114);
      gj_convTransposeB_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_sources/type_cast_2179/SplitProtocol/Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_sources/type_cast_2179/SplitProtocol/Sample/$exit
      -- 
    ra_5710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2179_inst_ack_0, ack => convTransposeB_CP_4753_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_sources/type_cast_2179/SplitProtocol/Update/ca
      -- CP-element group 117: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_sources/type_cast_2179/SplitProtocol/Update/$exit
      -- 
    ca_5715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2179_inst_ack_1, ack => convTransposeB_CP_4753_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	122 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_req
      -- CP-element group 118: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_sources/type_cast_2179/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_sources/type_cast_2179/$exit
      -- CP-element group 118: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2176/phi_stmt_2176_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2176/$exit
      -- 
    phi_stmt_2176_req_5716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2176_req_5716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(118), ack => phi_stmt_2176_req_0); -- 
    convTransposeB_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(116) & convTransposeB_CP_4753_elements(117);
      gj_convTransposeB_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	69 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2192/SplitProtocol/Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2192/SplitProtocol/Sample/$exit
      -- 
    ra_5733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2192_inst_ack_0, ack => convTransposeB_CP_4753_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	69 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2192/SplitProtocol/Update/ca
      -- CP-element group 120: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2192/SplitProtocol/Update/$exit
      -- 
    ca_5738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2192_inst_ack_1, ack => convTransposeB_CP_4753_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_req
      -- CP-element group 121: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2192/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/type_cast_2192/$exit
      -- CP-element group 121: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2189/phi_stmt_2189_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/phi_stmt_2189/$exit
      -- 
    phi_stmt_2189_req_5739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2189_req_5739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4753_elements(121), ack => phi_stmt_2189_req_0); -- 
    convTransposeB_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(119) & convTransposeB_CP_4753_elements(120);
      gj_convTransposeB_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: 	118 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1853/ifx_xthen_ifx_xend128_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(115) & convTransposeB_CP_4753_elements(118) & convTransposeB_CP_4753_elements(121);
      gj_convTransposeB_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	112 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_1853/merge_stmt_2175_PhiAck/$entry
      -- CP-element group 123: 	 branch_block_stmt_1853/merge_stmt_2175_PhiReqMerge
      -- 
    convTransposeB_CP_4753_elements(123) <= OrReduce(convTransposeB_CP_4753_elements(112) & convTransposeB_CP_4753_elements(122));
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1853/merge_stmt_2175_PhiAck/phi_stmt_2176_ack
      -- 
    phi_stmt_2176_ack_5744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2176_ack_0, ack => convTransposeB_CP_4753_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1853/merge_stmt_2175_PhiAck/phi_stmt_2183_ack
      -- 
    phi_stmt_2183_ack_5745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2183_ack_0, ack => convTransposeB_CP_4753_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1853/merge_stmt_2175_PhiAck/phi_stmt_2189_ack
      -- 
    phi_stmt_2189_ack_5746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2189_ack_0, ack => convTransposeB_CP_4753_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1853/merge_stmt_2175_PhiAck/$exit
      -- 
    convTransposeB_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4753_elements(124) & convTransposeB_CP_4753_elements(125) & convTransposeB_CP_4753_elements(126);
      gj_convTransposeB_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4753_elements(127), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom86_2095_resized : std_logic_vector(13 downto 0);
    signal R_idxprom86_2095_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2072_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2072_scaled : std_logic_vector(13 downto 0);
    signal add45_1927 : std_logic_vector(15 downto 0);
    signal add58_1938 : std_logic_vector(15 downto 0);
    signal add77_2048 : std_logic_vector(63 downto 0);
    signal add79_2058 : std_logic_vector(63 downto 0);
    signal add91_2112 : std_logic_vector(31 downto 0);
    signal add98_2130 : std_logic_vector(15 downto 0);
    signal add_1905 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2006 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2073_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2073_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2073_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2073_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2073_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2073_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2096_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2096_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2096_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2096_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2096_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2096_root_address : std_logic_vector(13 downto 0);
    signal arrayidx82_2075 : std_logic_vector(31 downto 0);
    signal arrayidx87_2098 : std_logic_vector(31 downto 0);
    signal call11_1874 : std_logic_vector(15 downto 0);
    signal call13_1877 : std_logic_vector(15 downto 0);
    signal call14_1880 : std_logic_vector(15 downto 0);
    signal call15_1883 : std_logic_vector(15 downto 0);
    signal call16_1896 : std_logic_vector(15 downto 0);
    signal call18_1908 : std_logic_vector(15 downto 0);
    signal call1_1859 : std_logic_vector(15 downto 0);
    signal call20_1911 : std_logic_vector(15 downto 0);
    signal call22_1914 : std_logic_vector(15 downto 0);
    signal call3_1862 : std_logic_vector(15 downto 0);
    signal call5_1865 : std_logic_vector(15 downto 0);
    signal call7_1868 : std_logic_vector(15 downto 0);
    signal call9_1871 : std_logic_vector(15 downto 0);
    signal call_1856 : std_logic_vector(15 downto 0);
    signal cmp106_2143 : std_logic_vector(0 downto 0);
    signal cmp117_2168 : std_logic_vector(0 downto 0);
    signal cmp_2117 : std_logic_vector(0 downto 0);
    signal conv112_2163 : std_logic_vector(31 downto 0);
    signal conv115_1959 : std_logic_vector(31 downto 0);
    signal conv17_1900 : std_logic_vector(31 downto 0);
    signal conv65_2030 : std_logic_vector(63 downto 0);
    signal conv68_1947 : std_logic_vector(63 downto 0);
    signal conv70_2034 : std_logic_vector(63 downto 0);
    signal conv73_1951 : std_logic_vector(63 downto 0);
    signal conv75_2038 : std_logic_vector(63 downto 0);
    signal conv90_2106 : std_logic_vector(31 downto 0);
    signal conv94_1955 : std_logic_vector(31 downto 0);
    signal conv_1887 : std_logic_vector(31 downto 0);
    signal idxprom86_2091 : std_logic_vector(63 downto 0);
    signal idxprom_2068 : std_logic_vector(63 downto 0);
    signal inc110_2147 : std_logic_vector(15 downto 0);
    signal inc110x_xinput_dim0x_x2_2152 : std_logic_vector(15 downto 0);
    signal inc_2138 : std_logic_vector(15 downto 0);
    signal indvar_1968 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2201 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2189 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1989 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2183 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1982 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2159 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2176 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1975 : std_logic_vector(15 downto 0);
    signal mul54_2021 : std_logic_vector(15 downto 0);
    signal mul76_2043 : std_logic_vector(63 downto 0);
    signal mul78_2053 : std_logic_vector(63 downto 0);
    signal mul_2011 : std_logic_vector(15 downto 0);
    signal ptr_deref_2078_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2078_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2078_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2078_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2078_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2100_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2100_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2100_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2100_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2100_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2100_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_1893 : std_logic_vector(31 downto 0);
    signal shr116132_1965 : std_logic_vector(31 downto 0);
    signal shr131_1921 : std_logic_vector(15 downto 0);
    signal shr81_2064 : std_logic_vector(31 downto 0);
    signal shr85_2085 : std_logic_vector(63 downto 0);
    signal sub48_2016 : std_logic_vector(15 downto 0);
    signal sub61_1943 : std_logic_vector(15 downto 0);
    signal sub62_2026 : std_logic_vector(15 downto 0);
    signal sub_1932 : std_logic_vector(15 downto 0);
    signal tmp1_2001 : std_logic_vector(31 downto 0);
    signal tmp83_2079 : std_logic_vector(63 downto 0);
    signal type_cast_1891_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1919_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1925_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1936_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1963_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1972_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1974_wire : std_logic_vector(31 downto 0);
    signal type_cast_1979_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1981_wire : std_logic_vector(15 downto 0);
    signal type_cast_1985_wire : std_logic_vector(15 downto 0);
    signal type_cast_1988_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1992_wire : std_logic_vector(15 downto 0);
    signal type_cast_1994_wire : std_logic_vector(15 downto 0);
    signal type_cast_1999_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2062_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2083_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2089_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2110_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2128_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2136_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2156_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2179_wire : std_logic_vector(15 downto 0);
    signal type_cast_2182_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2186_wire : std_logic_vector(15 downto 0);
    signal type_cast_2188_wire : std_logic_vector(15 downto 0);
    signal type_cast_2192_wire : std_logic_vector(15 downto 0);
    signal type_cast_2194_wire : std_logic_vector(15 downto 0);
    signal type_cast_2199_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2207_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2073_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2073_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2073_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2073_resized_base_address <= "00000000000000";
    array_obj_ref_2096_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2096_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2096_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2096_resized_base_address <= "00000000000000";
    ptr_deref_2078_word_offset_0 <= "00000000000000";
    ptr_deref_2100_word_offset_0 <= "00000000000000";
    type_cast_1891_wire_constant <= "00000000000000000000000000010000";
    type_cast_1919_wire_constant <= "0000000000000010";
    type_cast_1925_wire_constant <= "1111111111111111";
    type_cast_1936_wire_constant <= "1111111111111111";
    type_cast_1963_wire_constant <= "00000000000000000000000000000001";
    type_cast_1972_wire_constant <= "00000000000000000000000000000000";
    type_cast_1979_wire_constant <= "0000000000000000";
    type_cast_1988_wire_constant <= "0000000000000000";
    type_cast_1999_wire_constant <= "00000000000000000000000000000100";
    type_cast_2062_wire_constant <= "00000000000000000000000000000010";
    type_cast_2083_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2089_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2110_wire_constant <= "00000000000000000000000000000100";
    type_cast_2128_wire_constant <= "0000000000000100";
    type_cast_2136_wire_constant <= "0000000000000001";
    type_cast_2156_wire_constant <= "0000000000000000";
    type_cast_2182_wire_constant <= "0000000000000000";
    type_cast_2199_wire_constant <= "00000000000000000000000000000001";
    type_cast_2207_wire_constant <= "0000000000000001";
    phi_stmt_1968: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1972_wire_constant & type_cast_1974_wire;
      req <= phi_stmt_1968_req_0 & phi_stmt_1968_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1968",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1968_ack_0,
          idata => idata,
          odata => indvar_1968,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1968
    phi_stmt_1975: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1979_wire_constant & type_cast_1981_wire;
      req <= phi_stmt_1975_req_0 & phi_stmt_1975_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1975",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1975_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1975,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1975
    phi_stmt_1982: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1985_wire & type_cast_1988_wire_constant;
      req <= phi_stmt_1982_req_0 & phi_stmt_1982_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1982",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1982_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1982,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1982
    phi_stmt_1989: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1992_wire & type_cast_1994_wire;
      req <= phi_stmt_1989_req_0 & phi_stmt_1989_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1989",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1989_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1989,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1989
    phi_stmt_2176: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2179_wire & type_cast_2182_wire_constant;
      req <= phi_stmt_2176_req_0 & phi_stmt_2176_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2176",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2176_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2176,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2176
    phi_stmt_2183: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2186_wire & type_cast_2188_wire;
      req <= phi_stmt_2183_req_0 & phi_stmt_2183_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2183",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2183_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2183,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2183
    phi_stmt_2189: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2192_wire & type_cast_2194_wire;
      req <= phi_stmt_2189_req_0 & phi_stmt_2189_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2189",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2189_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2189,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2189
    -- flow-through select operator MUX_2158_inst
    input_dim1x_x2_2159 <= type_cast_2156_wire_constant when (cmp106_2143(0) /=  '0') else inc_2138;
    addr_of_2074_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2074_final_reg_req_0;
      addr_of_2074_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2074_final_reg_req_1;
      addr_of_2074_final_reg_ack_1<= rack(0);
      addr_of_2074_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2074_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2073_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_2075,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2097_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2097_final_reg_req_0;
      addr_of_2097_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2097_final_reg_req_1;
      addr_of_2097_final_reg_ack_1<= rack(0);
      addr_of_2097_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2097_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2096_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2098,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1886_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1886_inst_req_0;
      type_cast_1886_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1886_inst_req_1;
      type_cast_1886_inst_ack_1<= rack(0);
      type_cast_1886_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1886_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_1883,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1887,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1899_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1899_inst_req_0;
      type_cast_1899_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1899_inst_req_1;
      type_cast_1899_inst_ack_1<= rack(0);
      type_cast_1899_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1899_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1896,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1900,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1946_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1946_inst_req_0;
      type_cast_1946_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1946_inst_req_1;
      type_cast_1946_inst_ack_1<= rack(0);
      type_cast_1946_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1946_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_1914,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_1947,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1950_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1950_inst_req_0;
      type_cast_1950_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1950_inst_req_1;
      type_cast_1950_inst_ack_1<= rack(0);
      type_cast_1950_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1950_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_1911,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_1951,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1954_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1954_inst_req_0;
      type_cast_1954_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1954_inst_req_1;
      type_cast_1954_inst_ack_1<= rack(0);
      type_cast_1954_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1954_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_1862,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_1955,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1958_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1958_inst_req_0;
      type_cast_1958_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1958_inst_req_1;
      type_cast_1958_inst_ack_1<= rack(0);
      type_cast_1958_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1958_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1856,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_1959,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1974_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1974_inst_req_0;
      type_cast_1974_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1974_inst_req_1;
      type_cast_1974_inst_ack_1<= rack(0);
      type_cast_1974_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1974_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2201,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1974_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1981_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1981_inst_req_0;
      type_cast_1981_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1981_inst_req_1;
      type_cast_1981_inst_ack_1<= rack(0);
      type_cast_1981_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1981_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2176,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1981_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1985_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1985_inst_req_0;
      type_cast_1985_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1985_inst_req_1;
      type_cast_1985_inst_ack_1<= rack(0);
      type_cast_1985_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1985_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2183,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1985_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1992_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1992_inst_req_0;
      type_cast_1992_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1992_inst_req_1;
      type_cast_1992_inst_ack_1<= rack(0);
      type_cast_1992_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1992_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr131_1921,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1992_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1994_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1994_inst_req_0;
      type_cast_1994_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1994_inst_req_1;
      type_cast_1994_inst_ack_1<= rack(0);
      type_cast_1994_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1994_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2189,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1994_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2029_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2029_inst_req_0;
      type_cast_2029_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2029_inst_req_1;
      type_cast_2029_inst_ack_1<= rack(0);
      type_cast_2029_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2029_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1975,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2030,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2033_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2033_inst_req_0;
      type_cast_2033_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2033_inst_req_1;
      type_cast_2033_inst_ack_1<= rack(0);
      type_cast_2033_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2033_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_2026,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2034,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2037_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2037_inst_req_0;
      type_cast_2037_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2037_inst_req_1;
      type_cast_2037_inst_ack_1<= rack(0);
      type_cast_2037_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2037_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_2016,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2038,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2067_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2067_inst_req_0;
      type_cast_2067_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2067_inst_req_1;
      type_cast_2067_inst_ack_1<= rack(0);
      type_cast_2067_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2067_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr81_2064,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2068,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2105_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2105_inst_req_0;
      type_cast_2105_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2105_inst_req_1;
      type_cast_2105_inst_ack_1<= rack(0);
      type_cast_2105_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2105_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1975,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_2106,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2146_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2146_inst_req_0;
      type_cast_2146_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2146_inst_req_1;
      type_cast_2146_inst_ack_1<= rack(0);
      type_cast_2146_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2146_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp106_2143,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc110_2147,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2162_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2162_inst_req_0;
      type_cast_2162_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2162_inst_req_1;
      type_cast_2162_inst_ack_1<= rack(0);
      type_cast_2162_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2162_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2152,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2163,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2179_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2179_inst_req_0;
      type_cast_2179_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2179_inst_req_1;
      type_cast_2179_inst_ack_1<= rack(0);
      type_cast_2179_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2179_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add98_2130,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2179_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2186_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2186_inst_req_0;
      type_cast_2186_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2186_inst_req_1;
      type_cast_2186_inst_ack_1<= rack(0);
      type_cast_2186_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2186_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2159,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2186_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2188_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2188_inst_req_0;
      type_cast_2188_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2188_inst_req_1;
      type_cast_2188_inst_ack_1<= rack(0);
      type_cast_2188_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2188_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1982,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2188_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2192_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2192_inst_req_0;
      type_cast_2192_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2192_inst_req_1;
      type_cast_2192_inst_ack_1<= rack(0);
      type_cast_2192_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2192_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1989,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2192_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2194_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2194_inst_req_0;
      type_cast_2194_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2194_inst_req_1;
      type_cast_2194_inst_ack_1<= rack(0);
      type_cast_2194_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2194_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2152,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2194_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2073_index_1_rename
    process(R_idxprom_2072_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2072_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2072_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2073_index_1_resize
    process(idxprom_2068) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2068;
      ov := iv(13 downto 0);
      R_idxprom_2072_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2073_root_address_inst
    process(array_obj_ref_2073_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2073_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2073_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2096_index_1_rename
    process(R_idxprom86_2095_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom86_2095_resized;
      ov(13 downto 0) := iv;
      R_idxprom86_2095_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2096_index_1_resize
    process(idxprom86_2091) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom86_2091;
      ov := iv(13 downto 0);
      R_idxprom86_2095_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2096_root_address_inst
    process(array_obj_ref_2096_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2096_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2096_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2078_addr_0
    process(ptr_deref_2078_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2078_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2078_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2078_base_resize
    process(arrayidx82_2075) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_2075;
      ov := iv(13 downto 0);
      ptr_deref_2078_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2078_gather_scatter
    process(ptr_deref_2078_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2078_data_0;
      ov(63 downto 0) := iv;
      tmp83_2079 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2078_root_address_inst
    process(ptr_deref_2078_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2078_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2078_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2100_addr_0
    process(ptr_deref_2100_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2100_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2100_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2100_base_resize
    process(arrayidx87_2098) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2098;
      ov := iv(13 downto 0);
      ptr_deref_2100_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2100_gather_scatter
    process(tmp83_2079) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp83_2079;
      ov(63 downto 0) := iv;
      ptr_deref_2100_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2100_root_address_inst
    process(ptr_deref_2100_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2100_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2100_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2118_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2117;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2118_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2118_branch_req_0,
          ack0 => if_stmt_2118_branch_ack_0,
          ack1 => if_stmt_2118_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2169_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp117_2168;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2169_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2169_branch_req_0,
          ack0 => if_stmt_2169_branch_ack_0,
          ack1 => if_stmt_2169_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1926_inst
    process(call7_1868) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_1868, type_cast_1925_wire_constant, tmp_var);
      add45_1927 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1937_inst
    process(call9_1871) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_1871, type_cast_1936_wire_constant, tmp_var);
      add58_1938 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2015_inst
    process(sub_1932, mul_2011) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1932, mul_2011, tmp_var);
      sub48_2016 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2025_inst
    process(sub61_1943, mul54_2021) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_1943, mul54_2021, tmp_var);
      sub62_2026 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2129_inst
    process(input_dim2x_x1_1975) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1975, type_cast_2128_wire_constant, tmp_var);
      add98_2130 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2137_inst
    process(input_dim1x_x1_1982) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1982, type_cast_2136_wire_constant, tmp_var);
      inc_2138 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2151_inst
    process(inc110_2147, input_dim0x_x2_1989) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc110_2147, input_dim0x_x2_1989, tmp_var);
      inc110x_xinput_dim0x_x2_2152 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2005_inst
    process(add_1905, tmp1_2001) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_1905, tmp1_2001, tmp_var);
      add_src_0x_x0_2006 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2111_inst
    process(conv90_2106) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv90_2106, type_cast_2110_wire_constant, tmp_var);
      add91_2112 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2200_inst
    process(indvar_1968) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1968, type_cast_2199_wire_constant, tmp_var);
      indvarx_xnext_2201 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2047_inst
    process(mul76_2043, conv70_2034) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_2043, conv70_2034, tmp_var);
      add77_2048 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2057_inst
    process(mul78_2053, conv65_2030) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_2053, conv65_2030, tmp_var);
      add79_2058 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2090_inst
    process(shr85_2085) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr85_2085, type_cast_2089_wire_constant, tmp_var);
      idxprom86_2091 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2142_inst
    process(inc_2138, call1_1859) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2138, call1_1859, tmp_var);
      cmp106_2143 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2167_inst
    process(conv112_2163, shr116132_1965) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2163, shr116132_1965, tmp_var);
      cmp117_2168 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1920_inst
    process(call_1856) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1856, type_cast_1919_wire_constant, tmp_var);
      shr131_1921 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1964_inst
    process(conv115_1959) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_1959, type_cast_1963_wire_constant, tmp_var);
      shr116132_1965 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2063_inst
    process(add_src_0x_x0_2006) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2006, type_cast_2062_wire_constant, tmp_var);
      shr81_2064 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2084_inst
    process(add79_2058) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_2058, type_cast_2083_wire_constant, tmp_var);
      shr85_2085 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2010_inst
    process(input_dim0x_x2_1989, call13_1877) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_1989, call13_1877, tmp_var);
      mul_2011 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2020_inst
    process(input_dim1x_x1_1982, call13_1877) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_1982, call13_1877, tmp_var);
      mul54_2021 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2000_inst
    process(indvar_1968) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1968, type_cast_1999_wire_constant, tmp_var);
      tmp1_2001 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2042_inst
    process(conv75_2038, conv73_1951) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_2038, conv73_1951, tmp_var);
      mul76_2043 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2052_inst
    process(add77_2048, conv68_1947) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_2048, conv68_1947, tmp_var);
      mul78_2053 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1904_inst
    process(shl_1893, conv17_1900) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1893, conv17_1900, tmp_var);
      add_1905 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1892_inst
    process(conv_1887) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_1887, type_cast_1891_wire_constant, tmp_var);
      shl_1893 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1931_inst
    process(add45_1927, call14_1880) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_1927, call14_1880, tmp_var);
      sub_1932 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1942_inst
    process(add58_1938, call14_1880) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_1938, call14_1880, tmp_var);
      sub61_1943 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2116_inst
    process(add91_2112, conv94_1955) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add91_2112, conv94_1955, tmp_var);
      cmp_2117 <= tmp_var; --
    end process;
    -- shared split operator group (29) : array_obj_ref_2073_index_offset 
    ApIntAdd_group_29: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2072_scaled;
      array_obj_ref_2073_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2073_index_offset_req_0;
      array_obj_ref_2073_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2073_index_offset_req_1;
      array_obj_ref_2073_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_29_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : array_obj_ref_2096_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom86_2095_scaled;
      array_obj_ref_2096_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2096_index_offset_req_0;
      array_obj_ref_2096_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2096_index_offset_req_1;
      array_obj_ref_2096_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared load operator group (0) : ptr_deref_2078_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2078_load_0_req_0;
      ptr_deref_2078_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2078_load_0_req_1;
      ptr_deref_2078_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2078_word_address_0;
      ptr_deref_2078_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2100_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2100_store_0_req_0;
      ptr_deref_2100_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2100_store_0_req_1;
      ptr_deref_2100_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2100_word_address_0;
      data_in <= ptr_deref_2100_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1855_inst RPIPE_Block1_start_1861_inst RPIPE_Block1_start_1858_inst RPIPE_Block1_start_1913_inst RPIPE_Block1_start_1910_inst RPIPE_Block1_start_1907_inst RPIPE_Block1_start_1895_inst RPIPE_Block1_start_1882_inst RPIPE_Block1_start_1879_inst RPIPE_Block1_start_1876_inst RPIPE_Block1_start_1873_inst RPIPE_Block1_start_1870_inst RPIPE_Block1_start_1867_inst RPIPE_Block1_start_1864_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block1_start_1855_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block1_start_1861_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block1_start_1858_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_1913_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_1910_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_1907_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_1895_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_1882_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_1879_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_1876_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_1873_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_1870_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_1867_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_1864_inst_req_0;
      RPIPE_Block1_start_1855_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block1_start_1861_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block1_start_1858_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_1913_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_1910_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_1907_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_1895_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_1882_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_1879_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_1876_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_1873_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_1870_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_1867_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_1864_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block1_start_1855_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block1_start_1861_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block1_start_1858_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_1913_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_1910_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_1907_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_1895_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_1882_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_1879_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_1876_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_1873_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_1870_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_1867_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_1864_inst_req_1;
      RPIPE_Block1_start_1855_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block1_start_1861_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block1_start_1858_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_1913_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_1910_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_1907_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_1895_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_1882_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_1879_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_1876_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_1873_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_1870_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_1867_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_1864_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_1856 <= data_out(223 downto 208);
      call3_1862 <= data_out(207 downto 192);
      call1_1859 <= data_out(191 downto 176);
      call22_1914 <= data_out(175 downto 160);
      call20_1911 <= data_out(159 downto 144);
      call18_1908 <= data_out(143 downto 128);
      call16_1896 <= data_out(127 downto 112);
      call15_1883 <= data_out(111 downto 96);
      call14_1880 <= data_out(95 downto 80);
      call13_1877 <= data_out(79 downto 64);
      call11_1874 <= data_out(63 downto 48);
      call9_1871 <= data_out(47 downto 32);
      call7_1868 <= data_out(31 downto 16);
      call5_1865 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2205_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2205_inst_req_0;
      WPIPE_Block1_done_2205_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2205_inst_req_1;
      WPIPE_Block1_done_2205_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2207_wire_constant;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_5763_start: Boolean;
  signal convTransposeC_CP_5763_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block2_start_2234_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2243_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2271_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2228_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2234_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2243_inst_ack_1 : boolean;
  signal type_cast_2260_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2271_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2268_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2237_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2240_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2237_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2228_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2225_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2237_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2268_inst_req_0 : boolean;
  signal type_cast_2260_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2225_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2256_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2225_inst_ack_0 : boolean;
  signal type_cast_2247_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2231_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2231_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2225_inst_ack_1 : boolean;
  signal type_cast_2247_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2256_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2271_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2268_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2234_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2256_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2237_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2234_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2231_inst_req_1 : boolean;
  signal type_cast_2247_inst_req_1 : boolean;
  signal type_cast_2260_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2231_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2240_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2240_inst_ack_0 : boolean;
  signal type_cast_2247_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2271_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2240_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2256_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2243_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2228_inst_ack_0 : boolean;
  signal type_cast_2260_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2243_inst_ack_0 : boolean;
  signal type_cast_2311_inst_req_1 : boolean;
  signal type_cast_2319_inst_req_0 : boolean;
  signal type_cast_2319_inst_ack_0 : boolean;
  signal type_cast_2315_inst_req_1 : boolean;
  signal type_cast_2315_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2274_inst_ack_1 : boolean;
  signal type_cast_2315_inst_req_0 : boolean;
  signal type_cast_2315_inst_ack_0 : boolean;
  signal type_cast_2307_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2274_inst_req_1 : boolean;
  signal type_cast_2307_inst_req_1 : boolean;
  signal type_cast_2319_inst_req_1 : boolean;
  signal type_cast_2319_inst_ack_1 : boolean;
  signal type_cast_2311_inst_ack_1 : boolean;
  signal type_cast_2311_inst_ack_0 : boolean;
  signal type_cast_2311_inst_req_0 : boolean;
  signal type_cast_2307_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2274_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2228_inst_req_0 : boolean;
  signal type_cast_2307_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2274_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2222_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2268_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2216_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2216_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2216_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2216_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2219_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2219_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2219_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2219_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2222_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2222_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2222_inst_req_1 : boolean;
  signal type_cast_2401_inst_req_0 : boolean;
  signal type_cast_2401_inst_ack_0 : boolean;
  signal type_cast_2401_inst_req_1 : boolean;
  signal type_cast_2401_inst_ack_1 : boolean;
  signal type_cast_2405_inst_req_0 : boolean;
  signal type_cast_2405_inst_ack_0 : boolean;
  signal type_cast_2405_inst_req_1 : boolean;
  signal type_cast_2405_inst_ack_1 : boolean;
  signal type_cast_2409_inst_req_0 : boolean;
  signal type_cast_2409_inst_ack_0 : boolean;
  signal type_cast_2409_inst_req_1 : boolean;
  signal type_cast_2409_inst_ack_1 : boolean;
  signal type_cast_2439_inst_req_0 : boolean;
  signal type_cast_2439_inst_ack_0 : boolean;
  signal type_cast_2439_inst_req_1 : boolean;
  signal type_cast_2439_inst_ack_1 : boolean;
  signal array_obj_ref_2445_index_offset_req_0 : boolean;
  signal array_obj_ref_2445_index_offset_ack_0 : boolean;
  signal array_obj_ref_2445_index_offset_req_1 : boolean;
  signal array_obj_ref_2445_index_offset_ack_1 : boolean;
  signal addr_of_2446_final_reg_req_0 : boolean;
  signal addr_of_2446_final_reg_ack_0 : boolean;
  signal addr_of_2446_final_reg_req_1 : boolean;
  signal addr_of_2446_final_reg_ack_1 : boolean;
  signal ptr_deref_2450_load_0_req_0 : boolean;
  signal ptr_deref_2450_load_0_ack_0 : boolean;
  signal ptr_deref_2450_load_0_req_1 : boolean;
  signal ptr_deref_2450_load_0_ack_1 : boolean;
  signal array_obj_ref_2468_index_offset_req_0 : boolean;
  signal array_obj_ref_2468_index_offset_ack_0 : boolean;
  signal array_obj_ref_2468_index_offset_req_1 : boolean;
  signal array_obj_ref_2468_index_offset_ack_1 : boolean;
  signal addr_of_2469_final_reg_req_0 : boolean;
  signal addr_of_2469_final_reg_ack_0 : boolean;
  signal addr_of_2469_final_reg_req_1 : boolean;
  signal addr_of_2469_final_reg_ack_1 : boolean;
  signal ptr_deref_2472_store_0_req_0 : boolean;
  signal ptr_deref_2472_store_0_ack_0 : boolean;
  signal ptr_deref_2472_store_0_req_1 : boolean;
  signal ptr_deref_2472_store_0_ack_1 : boolean;
  signal type_cast_2477_inst_req_0 : boolean;
  signal type_cast_2477_inst_ack_0 : boolean;
  signal type_cast_2477_inst_req_1 : boolean;
  signal type_cast_2477_inst_ack_1 : boolean;
  signal if_stmt_2490_branch_req_0 : boolean;
  signal if_stmt_2490_branch_ack_1 : boolean;
  signal if_stmt_2490_branch_ack_0 : boolean;
  signal type_cast_2518_inst_req_0 : boolean;
  signal type_cast_2518_inst_ack_0 : boolean;
  signal type_cast_2518_inst_req_1 : boolean;
  signal type_cast_2518_inst_ack_1 : boolean;
  signal type_cast_2534_inst_req_0 : boolean;
  signal type_cast_2534_inst_ack_0 : boolean;
  signal type_cast_2534_inst_req_1 : boolean;
  signal type_cast_2534_inst_ack_1 : boolean;
  signal if_stmt_2541_branch_req_0 : boolean;
  signal if_stmt_2541_branch_ack_1 : boolean;
  signal if_stmt_2541_branch_ack_0 : boolean;
  signal WPIPE_Block2_done_2577_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2577_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2577_inst_req_1 : boolean;
  signal WPIPE_Block2_done_2577_inst_ack_1 : boolean;
  signal phi_stmt_2340_req_0 : boolean;
  signal phi_stmt_2347_req_1 : boolean;
  signal phi_stmt_2354_req_1 : boolean;
  signal type_cast_2366_inst_req_0 : boolean;
  signal type_cast_2366_inst_ack_0 : boolean;
  signal type_cast_2366_inst_req_1 : boolean;
  signal type_cast_2366_inst_ack_1 : boolean;
  signal phi_stmt_2361_req_1 : boolean;
  signal type_cast_2346_inst_req_0 : boolean;
  signal type_cast_2346_inst_ack_0 : boolean;
  signal type_cast_2346_inst_req_1 : boolean;
  signal type_cast_2346_inst_ack_1 : boolean;
  signal phi_stmt_2340_req_1 : boolean;
  signal type_cast_2350_inst_req_0 : boolean;
  signal type_cast_2350_inst_ack_0 : boolean;
  signal type_cast_2350_inst_req_1 : boolean;
  signal type_cast_2350_inst_ack_1 : boolean;
  signal phi_stmt_2347_req_0 : boolean;
  signal type_cast_2357_inst_req_0 : boolean;
  signal type_cast_2357_inst_ack_0 : boolean;
  signal type_cast_2357_inst_req_1 : boolean;
  signal type_cast_2357_inst_ack_1 : boolean;
  signal phi_stmt_2354_req_0 : boolean;
  signal type_cast_2364_inst_req_0 : boolean;
  signal type_cast_2364_inst_ack_0 : boolean;
  signal type_cast_2364_inst_req_1 : boolean;
  signal type_cast_2364_inst_ack_1 : boolean;
  signal phi_stmt_2361_req_0 : boolean;
  signal phi_stmt_2340_ack_0 : boolean;
  signal phi_stmt_2347_ack_0 : boolean;
  signal phi_stmt_2354_ack_0 : boolean;
  signal phi_stmt_2361_ack_0 : boolean;
  signal phi_stmt_2548_req_1 : boolean;
  signal type_cast_2558_inst_req_0 : boolean;
  signal type_cast_2558_inst_ack_0 : boolean;
  signal type_cast_2558_inst_req_1 : boolean;
  signal type_cast_2558_inst_ack_1 : boolean;
  signal phi_stmt_2555_req_0 : boolean;
  signal type_cast_2564_inst_req_0 : boolean;
  signal type_cast_2564_inst_ack_0 : boolean;
  signal type_cast_2564_inst_req_1 : boolean;
  signal type_cast_2564_inst_ack_1 : boolean;
  signal phi_stmt_2561_req_0 : boolean;
  signal type_cast_2551_inst_req_0 : boolean;
  signal type_cast_2551_inst_ack_0 : boolean;
  signal type_cast_2551_inst_req_1 : boolean;
  signal type_cast_2551_inst_ack_1 : boolean;
  signal phi_stmt_2548_req_0 : boolean;
  signal type_cast_2560_inst_req_0 : boolean;
  signal type_cast_2560_inst_ack_0 : boolean;
  signal type_cast_2560_inst_req_1 : boolean;
  signal type_cast_2560_inst_ack_1 : boolean;
  signal phi_stmt_2555_req_1 : boolean;
  signal type_cast_2566_inst_req_0 : boolean;
  signal type_cast_2566_inst_ack_0 : boolean;
  signal type_cast_2566_inst_req_1 : boolean;
  signal type_cast_2566_inst_ack_1 : boolean;
  signal phi_stmt_2561_req_1 : boolean;
  signal phi_stmt_2548_ack_0 : boolean;
  signal phi_stmt_2555_ack_0 : boolean;
  signal phi_stmt_2561_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_5763_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5763_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_5763_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5763_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_5763: Block -- control-path 
    signal convTransposeC_CP_5763_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_5763_elements(0) <= convTransposeC_CP_5763_start;
    convTransposeC_CP_5763_symbol <= convTransposeC_CP_5763_elements(78);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2260_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2247_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2260_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2247_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2260_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2247_Update/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2214/$entry
      -- CP-element group 0: 	 branch_block_stmt_2214/branch_block_stmt_2214__entry__
      -- CP-element group 0: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275__entry__
      -- CP-element group 0: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/$entry
      -- CP-element group 0: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2216_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2216_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2216_Sample/rr
      -- 
    cr_5984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(0), ack => type_cast_2260_inst_req_1); -- 
    cr_5956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(0), ack => type_cast_2247_inst_req_1); -- 
    rr_5811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(0), ack => RPIPE_Block2_start_2216_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	87 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	90 
    -- CP-element group 1: 	92 
    -- CP-element group 1: 	93 
    -- CP-element group 1: 	95 
    -- CP-element group 1: 	96 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2214/merge_stmt_2547__exit__
      -- CP-element group 1: 	 branch_block_stmt_2214/assign_stmt_2573__entry__
      -- CP-element group 1: 	 branch_block_stmt_2214/assign_stmt_2573__exit__
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2214/assign_stmt_2573/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/assign_stmt_2573/$exit
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2340/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_sources/type_cast_2346/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_sources/type_cast_2346/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_sources/type_cast_2346/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_sources/type_cast_2346/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_sources/type_cast_2346/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_sources/type_cast_2346/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2347/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_sources/type_cast_2350/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_sources/type_cast_2350/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_sources/type_cast_2350/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_sources/type_cast_2350/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_sources/type_cast_2350/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_sources/type_cast_2350/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2354/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_sources/type_cast_2357/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_sources/type_cast_2357/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_sources/type_cast_2357/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_sources/type_cast_2357/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_sources/type_cast_2357/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_sources/type_cast_2357/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2361/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2364/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2364/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2364/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2364/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2364/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2364/SplitProtocol/Update/cr
      -- 
    rr_6512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(1), ack => type_cast_2346_inst_req_0); -- 
    cr_6517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(1), ack => type_cast_2346_inst_req_1); -- 
    rr_6535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(1), ack => type_cast_2350_inst_req_0); -- 
    cr_6540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(1), ack => type_cast_2350_inst_req_1); -- 
    rr_6558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(1), ack => type_cast_2357_inst_req_0); -- 
    cr_6563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(1), ack => type_cast_2357_inst_req_1); -- 
    rr_6581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(1), ack => type_cast_2364_inst_req_0); -- 
    cr_6586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(1), ack => type_cast_2364_inst_req_1); -- 
    convTransposeC_CP_5763_elements(1) <= convTransposeC_CP_5763_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2216_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2216_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2216_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2216_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2216_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2216_Update/cr
      -- 
    ra_5812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2216_inst_ack_0, ack => convTransposeC_CP_5763_elements(2)); -- 
    cr_5816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(2), ack => RPIPE_Block2_start_2216_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2216_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2216_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2216_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2219_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2219_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2219_Sample/rr
      -- 
    ca_5817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2216_inst_ack_1, ack => convTransposeC_CP_5763_elements(3)); -- 
    rr_5825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(3), ack => RPIPE_Block2_start_2219_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2219_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2219_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2219_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2219_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2219_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2219_Update/cr
      -- 
    ra_5826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2219_inst_ack_0, ack => convTransposeC_CP_5763_elements(4)); -- 
    cr_5830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(4), ack => RPIPE_Block2_start_2219_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2219_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2219_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2219_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2222_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2222_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2222_Sample/rr
      -- 
    ca_5831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2219_inst_ack_1, ack => convTransposeC_CP_5763_elements(5)); -- 
    rr_5839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(5), ack => RPIPE_Block2_start_2222_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2222_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2222_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2222_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2222_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2222_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2222_Update/cr
      -- 
    ra_5840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2222_inst_ack_0, ack => convTransposeC_CP_5763_elements(6)); -- 
    cr_5844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(6), ack => RPIPE_Block2_start_2222_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2225_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2225_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2225_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2222_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2222_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2222_Update/$exit
      -- 
    ca_5845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2222_inst_ack_1, ack => convTransposeC_CP_5763_elements(7)); -- 
    rr_5853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(7), ack => RPIPE_Block2_start_2225_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2225_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2225_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2225_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2225_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2225_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2225_Update/$entry
      -- 
    ra_5854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2225_inst_ack_0, ack => convTransposeC_CP_5763_elements(8)); -- 
    cr_5858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(8), ack => RPIPE_Block2_start_2225_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2225_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2225_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2228_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2225_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2228_Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2228_Sample/$entry
      -- 
    ca_5859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2225_inst_ack_1, ack => convTransposeC_CP_5763_elements(9)); -- 
    rr_5867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(9), ack => RPIPE_Block2_start_2228_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2228_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2228_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2228_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2228_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2228_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2228_update_start_
      -- 
    ra_5868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2228_inst_ack_0, ack => convTransposeC_CP_5763_elements(10)); -- 
    cr_5872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(10), ack => RPIPE_Block2_start_2228_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2228_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2231_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2231_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2231_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2228_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2228_update_completed_
      -- 
    ca_5873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2228_inst_ack_1, ack => convTransposeC_CP_5763_elements(11)); -- 
    rr_5881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(11), ack => RPIPE_Block2_start_2231_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2231_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2231_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2231_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2231_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2231_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2231_Update/cr
      -- 
    ra_5882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2231_inst_ack_0, ack => convTransposeC_CP_5763_elements(12)); -- 
    cr_5886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(12), ack => RPIPE_Block2_start_2231_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2234_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2231_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2231_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2234_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2231_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2234_sample_start_
      -- 
    ca_5887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2231_inst_ack_1, ack => convTransposeC_CP_5763_elements(13)); -- 
    rr_5895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(13), ack => RPIPE_Block2_start_2234_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2234_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2234_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2234_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2234_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2234_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2234_update_start_
      -- 
    ra_5896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2234_inst_ack_0, ack => convTransposeC_CP_5763_elements(14)); -- 
    cr_5900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(14), ack => RPIPE_Block2_start_2234_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2234_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2237_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2234_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2234_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2237_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2237_sample_start_
      -- 
    ca_5901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2234_inst_ack_1, ack => convTransposeC_CP_5763_elements(15)); -- 
    rr_5909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(15), ack => RPIPE_Block2_start_2237_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2237_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2237_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2237_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2237_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2237_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2237_sample_completed_
      -- 
    ra_5910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2237_inst_ack_0, ack => convTransposeC_CP_5763_elements(16)); -- 
    cr_5914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(16), ack => RPIPE_Block2_start_2237_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2237_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2237_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2237_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2240_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2240_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2240_Sample/rr
      -- 
    ca_5915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2237_inst_ack_1, ack => convTransposeC_CP_5763_elements(17)); -- 
    rr_5923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(17), ack => RPIPE_Block2_start_2240_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2240_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2240_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2240_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2240_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2240_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2240_Update/cr
      -- 
    ra_5924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2240_inst_ack_0, ack => convTransposeC_CP_5763_elements(18)); -- 
    cr_5928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(18), ack => RPIPE_Block2_start_2240_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2243_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2240_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2240_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2240_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2243_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2243_sample_start_
      -- 
    ca_5929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2240_inst_ack_1, ack => convTransposeC_CP_5763_elements(19)); -- 
    rr_5937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(19), ack => RPIPE_Block2_start_2243_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2243_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2243_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2243_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2243_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2243_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2243_Sample/ra
      -- 
    ra_5938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2243_inst_ack_0, ack => convTransposeC_CP_5763_elements(20)); -- 
    cr_5942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(20), ack => RPIPE_Block2_start_2243_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2243_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2243_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2243_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2247_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2247_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2247_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2256_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2256_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2256_Sample/$entry
      -- 
    ca_5943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2243_inst_ack_1, ack => convTransposeC_CP_5763_elements(21)); -- 
    rr_5951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(21), ack => type_cast_2247_inst_req_0); -- 
    rr_5965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(21), ack => RPIPE_Block2_start_2256_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2247_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2247_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2247_Sample/ra
      -- 
    ra_5952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2247_inst_ack_0, ack => convTransposeC_CP_5763_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2247_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2247_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2247_Update/ca
      -- 
    ca_5957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2247_inst_ack_1, ack => convTransposeC_CP_5763_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2256_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2256_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2256_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2256_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2256_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2256_Sample/$exit
      -- 
    ra_5966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2256_inst_ack_0, ack => convTransposeC_CP_5763_elements(24)); -- 
    cr_5970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(24), ack => RPIPE_Block2_start_2256_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2268_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2260_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2256_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2268_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2256_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2268_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2260_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2256_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2260_Sample/rr
      -- 
    ca_5971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2256_inst_ack_1, ack => convTransposeC_CP_5763_elements(25)); -- 
    rr_5979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(25), ack => type_cast_2260_inst_req_0); -- 
    rr_5993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(25), ack => RPIPE_Block2_start_2268_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2260_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2260_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2260_Sample/ra
      -- 
    ra_5980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2260_inst_ack_0, ack => convTransposeC_CP_5763_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2260_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2260_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/type_cast_2260_Update/$exit
      -- 
    ca_5985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2260_inst_ack_1, ack => convTransposeC_CP_5763_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2268_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2268_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2268_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2268_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2268_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2268_Update/$entry
      -- 
    ra_5994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2268_inst_ack_0, ack => convTransposeC_CP_5763_elements(28)); -- 
    cr_5998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(28), ack => RPIPE_Block2_start_2268_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2268_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2271_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2271_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2268_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2271_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2268_Update/ca
      -- 
    ca_5999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2268_inst_ack_1, ack => convTransposeC_CP_5763_elements(29)); -- 
    rr_6007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(29), ack => RPIPE_Block2_start_2271_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2271_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2271_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2271_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2271_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2271_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2271_sample_completed_
      -- 
    ra_6008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2271_inst_ack_0, ack => convTransposeC_CP_5763_elements(30)); -- 
    cr_6012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(30), ack => RPIPE_Block2_start_2271_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2271_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2271_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2274_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2274_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2271_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2274_Sample/rr
      -- 
    ca_6013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2271_inst_ack_1, ack => convTransposeC_CP_5763_elements(31)); -- 
    rr_6021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(31), ack => RPIPE_Block2_start_2274_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2274_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2274_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2274_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2274_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2274_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2274_Sample/$exit
      -- 
    ra_6022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2274_inst_ack_0, ack => convTransposeC_CP_5763_elements(32)); -- 
    cr_6026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(32), ack => RPIPE_Block2_start_2274_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2274_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2274_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/RPIPE_Block2_start_2274_Update/$exit
      -- 
    ca_6027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2274_inst_ack_1, ack => convTransposeC_CP_5763_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34: 	41 
    -- CP-element group 34: 	42 
    -- CP-element group 34:  members (28) 
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2311_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2307_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2307_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2311_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2311_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2319_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2319_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2311_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/$entry
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2319_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2319_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2315_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2311_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2315_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2315_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2315_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2307_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2319_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2319_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2307_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2311_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2315_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2315_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2307_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2307_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275__exit__
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337__entry__
      -- CP-element group 34: 	 branch_block_stmt_2214/assign_stmt_2217_to_assign_stmt_2275/$exit
      -- 
    cr_6057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(34), ack => type_cast_2311_inst_req_1); -- 
    rr_6080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(34), ack => type_cast_2319_inst_req_0); -- 
    cr_6071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(34), ack => type_cast_2315_inst_req_1); -- 
    rr_6066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(34), ack => type_cast_2315_inst_req_0); -- 
    cr_6043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(34), ack => type_cast_2307_inst_req_1); -- 
    cr_6085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(34), ack => type_cast_2319_inst_req_1); -- 
    rr_6052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(34), ack => type_cast_2311_inst_req_0); -- 
    rr_6038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(34), ack => type_cast_2307_inst_req_0); -- 
    convTransposeC_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(23) & convTransposeC_CP_5763_elements(27) & convTransposeC_CP_5763_elements(33);
      gj_convTransposeC_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2307_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2307_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2307_Sample/$exit
      -- 
    ra_6039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2307_inst_ack_0, ack => convTransposeC_CP_5763_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	43 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2307_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2307_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2307_Update/$exit
      -- 
    ca_6044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2307_inst_ack_1, ack => convTransposeC_CP_5763_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2311_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2311_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2311_Sample/$exit
      -- 
    ra_6053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2311_inst_ack_0, ack => convTransposeC_CP_5763_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	43 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2311_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2311_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2311_Update/ca
      -- 
    ca_6058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2311_inst_ack_1, ack => convTransposeC_CP_5763_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2315_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2315_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2315_sample_completed_
      -- 
    ra_6067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2315_inst_ack_0, ack => convTransposeC_CP_5763_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2315_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2315_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2315_update_completed_
      -- 
    ca_6072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2315_inst_ack_1, ack => convTransposeC_CP_5763_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2319_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2319_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2319_sample_completed_
      -- 
    ra_6081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2319_inst_ack_0, ack => convTransposeC_CP_5763_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	34 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2319_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2319_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/type_cast_2319_Update/ca
      -- 
    ca_6086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2319_inst_ack_1, ack => convTransposeC_CP_5763_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  place  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	36 
    -- CP-element group 43: 	38 
    -- CP-element group 43: 	40 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	79 
    -- CP-element group 43: 	80 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	82 
    -- CP-element group 43: 	83 
    -- CP-element group 43:  members (18) 
      -- CP-element group 43: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337/$exit
      -- CP-element group 43: 	 branch_block_stmt_2214/assign_stmt_2282_to_assign_stmt_2337__exit__
      -- CP-element group 43: 	 branch_block_stmt_2214/entry_whilex_xbody
      -- CP-element group 43: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2340/$entry
      -- CP-element group 43: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2347/$entry
      -- CP-element group 43: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2354/$entry
      -- CP-element group 43: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2361/$entry
      -- CP-element group 43: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/$entry
      -- CP-element group 43: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2366/$entry
      -- CP-element group 43: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2366/SplitProtocol/$entry
      -- CP-element group 43: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2366/SplitProtocol/Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2366/SplitProtocol/Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2366/SplitProtocol/Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2366/SplitProtocol/Update/cr
      -- 
    rr_6486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(43), ack => type_cast_2366_inst_req_0); -- 
    cr_6491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(43), ack => type_cast_2366_inst_req_1); -- 
    convTransposeC_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(36) & convTransposeC_CP_5763_elements(38) & convTransposeC_CP_5763_elements(40) & convTransposeC_CP_5763_elements(42);
      gj_convTransposeC_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	104 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2401_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2401_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2401_Sample/ra
      -- 
    ra_6098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2401_inst_ack_0, ack => convTransposeC_CP_5763_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	104 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	58 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2401_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2401_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2401_Update/ca
      -- 
    ca_6103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2401_inst_ack_1, ack => convTransposeC_CP_5763_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	104 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2405_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2405_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2405_Sample/ra
      -- 
    ra_6112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2405_inst_ack_0, ack => convTransposeC_CP_5763_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	104 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	58 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2405_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2405_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2405_Update/ca
      -- 
    ca_6117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2405_inst_ack_1, ack => convTransposeC_CP_5763_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	104 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2409_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2409_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2409_Sample/ra
      -- 
    ra_6126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2409_inst_ack_0, ack => convTransposeC_CP_5763_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	104 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2409_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2409_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2409_Update/ca
      -- 
    ca_6131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2409_inst_ack_1, ack => convTransposeC_CP_5763_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	104 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2439_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2439_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2439_Sample/ra
      -- 
    ra_6140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2439_inst_ack_0, ack => convTransposeC_CP_5763_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	104 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (16) 
      -- CP-element group 51: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2439_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2439_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2439_Update/ca
      -- CP-element group 51: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_index_resized_1
      -- CP-element group 51: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_index_scaled_1
      -- CP-element group 51: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_index_computed_1
      -- CP-element group 51: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_index_resize_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_index_resize_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_index_resize_1/index_resize_req
      -- CP-element group 51: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_index_resize_1/index_resize_ack
      -- CP-element group 51: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_index_scale_1/$entry
      -- CP-element group 51: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_index_scale_1/$exit
      -- CP-element group 51: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_index_scale_1/scale_rename_req
      -- CP-element group 51: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_index_scale_1/scale_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_final_index_sum_regn_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_final_index_sum_regn_Sample/req
      -- 
    ca_6145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2439_inst_ack_1, ack => convTransposeC_CP_5763_elements(51)); -- 
    req_6170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(51), ack => array_obj_ref_2445_index_offset_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	68 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_final_index_sum_regn_sample_complete
      -- CP-element group 52: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_final_index_sum_regn_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_final_index_sum_regn_Sample/ack
      -- 
    ack_6171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2445_index_offset_ack_0, ack => convTransposeC_CP_5763_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	104 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (11) 
      -- CP-element group 53: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2446_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_offset_calculated
      -- CP-element group 53: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_final_index_sum_regn_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_final_index_sum_regn_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2446_request/$entry
      -- CP-element group 53: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2446_request/req
      -- 
    ack_6176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2445_index_offset_ack_1, ack => convTransposeC_CP_5763_elements(53)); -- 
    req_6185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(53), ack => addr_of_2446_final_reg_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2446_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2446_request/$exit
      -- CP-element group 54: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2446_request/ack
      -- 
    ack_6186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2446_final_reg_ack_0, ack => convTransposeC_CP_5763_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	104 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (24) 
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2446_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2446_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2446_complete/ack
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_base_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_word_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_root_address_calculated
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_base_address_resized
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_base_addr_resize/$entry
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_base_addr_resize/$exit
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_base_addr_resize/base_resize_req
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_base_addr_resize/base_resize_ack
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_base_plus_offset/$entry
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_base_plus_offset/$exit
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_base_plus_offset/sum_rename_req
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_base_plus_offset/sum_rename_ack
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_word_addrgen/$entry
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_word_addrgen/$exit
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_word_addrgen/root_register_req
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_word_addrgen/root_register_ack
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Sample/word_access_start/word_0/rr
      -- 
    ack_6191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2446_final_reg_ack_1, ack => convTransposeC_CP_5763_elements(55)); -- 
    rr_6224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(55), ack => ptr_deref_2450_load_0_req_0); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Sample/word_access_start/word_0/ra
      -- 
    ra_6225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2450_load_0_ack_0, ack => convTransposeC_CP_5763_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	104 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Update/word_access_complete/word_0/ca
      -- CP-element group 57: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Update/ptr_deref_2450_Merge/$entry
      -- CP-element group 57: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Update/ptr_deref_2450_Merge/$exit
      -- CP-element group 57: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Update/ptr_deref_2450_Merge/merge_req
      -- CP-element group 57: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Update/ptr_deref_2450_Merge/merge_ack
      -- 
    ca_6236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2450_load_0_ack_1, ack => convTransposeC_CP_5763_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	47 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_final_index_sum_regn_Sample/req
      -- 
    req_6266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(58), ack => array_obj_ref_2468_index_offset_req_0); -- 
    convTransposeC_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(45) & convTransposeC_CP_5763_elements(47) & convTransposeC_CP_5763_elements(49);
      gj_convTransposeC_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	68 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_final_index_sum_regn_Sample/ack
      -- 
    ack_6267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2468_index_offset_ack_0, ack => convTransposeC_CP_5763_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	104 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2469_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2469_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2469_request/req
      -- 
    ack_6272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2468_index_offset_ack_1, ack => convTransposeC_CP_5763_elements(60)); -- 
    req_6281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(60), ack => addr_of_2469_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2469_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2469_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2469_request/ack
      -- 
    ack_6282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2469_final_reg_ack_0, ack => convTransposeC_CP_5763_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	104 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2469_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2469_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2469_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_word_addrgen/root_register_ack
      -- 
    ack_6287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2469_final_reg_ack_1, ack => convTransposeC_CP_5763_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Sample/ptr_deref_2472_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Sample/ptr_deref_2472_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Sample/ptr_deref_2472_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Sample/ptr_deref_2472_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Sample/word_access_start/word_0/rr
      -- 
    rr_6325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(63), ack => ptr_deref_2472_store_0_req_0); -- 
    convTransposeC_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(57) & convTransposeC_CP_5763_elements(62);
      gj_convTransposeC_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Sample/word_access_start/word_0/ra
      -- 
    ra_6326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2472_store_0_ack_0, ack => convTransposeC_CP_5763_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	104 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Update/word_access_complete/word_0/ca
      -- 
    ca_6337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2472_store_0_ack_1, ack => convTransposeC_CP_5763_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	104 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2477_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2477_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2477_Sample/ra
      -- 
    ra_6346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2477_inst_ack_0, ack => convTransposeC_CP_5763_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	104 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2477_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2477_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2477_Update/ca
      -- 
    ca_6351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2477_inst_ack_1, ack => convTransposeC_CP_5763_elements(67)); -- 
    -- CP-element group 68:  branch  join  transition  place  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	52 
    -- CP-element group 68: 	59 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (10) 
      -- CP-element group 68: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/$exit
      -- CP-element group 68: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489__exit__
      -- CP-element group 68: 	 branch_block_stmt_2214/if_stmt_2490__entry__
      -- CP-element group 68: 	 branch_block_stmt_2214/if_stmt_2490_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2214/if_stmt_2490_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_2214/if_stmt_2490_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_2214/if_stmt_2490_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_2214/R_cmp_2491_place
      -- CP-element group 68: 	 branch_block_stmt_2214/if_stmt_2490_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_2214/if_stmt_2490_else_link/$entry
      -- 
    branch_req_6359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(68), ack => if_stmt_2490_branch_req_0); -- 
    convTransposeC_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(52) & convTransposeC_CP_5763_elements(59) & convTransposeC_CP_5763_elements(65) & convTransposeC_CP_5763_elements(67);
      gj_convTransposeC_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	113 
    -- CP-element group 69: 	114 
    -- CP-element group 69: 	116 
    -- CP-element group 69: 	117 
    -- CP-element group 69: 	119 
    -- CP-element group 69: 	120 
    -- CP-element group 69:  members (40) 
      -- CP-element group 69: 	 branch_block_stmt_2214/merge_stmt_2496__exit__
      -- CP-element group 69: 	 branch_block_stmt_2214/assign_stmt_2502__entry__
      -- CP-element group 69: 	 branch_block_stmt_2214/assign_stmt_2502__exit__
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133
      -- CP-element group 69: 	 branch_block_stmt_2214/if_stmt_2490_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_2214/if_stmt_2490_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_2214/whilex_xbody_ifx_xthen
      -- CP-element group 69: 	 branch_block_stmt_2214/assign_stmt_2502/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/assign_stmt_2502/$exit
      -- CP-element group 69: 	 branch_block_stmt_2214/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_2214/merge_stmt_2496_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_2214/merge_stmt_2496_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/merge_stmt_2496_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_2214/merge_stmt_2496_PhiAck/dummy
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2548/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_sources/type_cast_2551/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_sources/type_cast_2551/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_sources/type_cast_2551/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_sources/type_cast_2551/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_sources/type_cast_2551/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_sources/type_cast_2551/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/Update/cr
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2561/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2566/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2566/SplitProtocol/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2566/SplitProtocol/Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2566/SplitProtocol/Sample/rr
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2566/SplitProtocol/Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2566/SplitProtocol/Update/cr
      -- 
    if_choice_transition_6364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2490_branch_ack_1, ack => convTransposeC_CP_5763_elements(69)); -- 
    rr_6696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(69), ack => type_cast_2551_inst_req_0); -- 
    cr_6701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(69), ack => type_cast_2551_inst_req_1); -- 
    rr_6719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(69), ack => type_cast_2560_inst_req_0); -- 
    cr_6724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(69), ack => type_cast_2560_inst_req_1); -- 
    rr_6742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(69), ack => type_cast_2566_inst_req_0); -- 
    cr_6747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(69), ack => type_cast_2566_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70: 	74 
    -- CP-element group 70:  members (21) 
      -- CP-element group 70: 	 branch_block_stmt_2214/merge_stmt_2504__exit__
      -- CP-element group 70: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540__entry__
      -- CP-element group 70: 	 branch_block_stmt_2214/if_stmt_2490_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_2214/if_stmt_2490_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_2214/whilex_xbody_ifx_xelse
      -- CP-element group 70: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/$entry
      -- CP-element group 70: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2518_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2518_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2518_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2518_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2518_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2518_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2534_update_start_
      -- CP-element group 70: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2534_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2534_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_2214/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_2214/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_2214/merge_stmt_2504_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_2214/merge_stmt_2504_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_2214/merge_stmt_2504_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_2214/merge_stmt_2504_PhiAck/dummy
      -- 
    else_choice_transition_6368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2490_branch_ack_0, ack => convTransposeC_CP_5763_elements(70)); -- 
    rr_6384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(70), ack => type_cast_2518_inst_req_0); -- 
    cr_6389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(70), ack => type_cast_2518_inst_req_1); -- 
    cr_6403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(70), ack => type_cast_2534_inst_req_1); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2518_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2518_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2518_Sample/ra
      -- 
    ra_6385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2518_inst_ack_0, ack => convTransposeC_CP_5763_elements(71)); -- 
    -- CP-element group 72:  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (6) 
      -- CP-element group 72: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2518_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2518_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2518_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2534_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2534_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2534_Sample/rr
      -- 
    ca_6390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2518_inst_ack_1, ack => convTransposeC_CP_5763_elements(72)); -- 
    rr_6398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(72), ack => type_cast_2534_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2534_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2534_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2534_Sample/ra
      -- 
    ra_6399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2534_inst_ack_0, ack => convTransposeC_CP_5763_elements(73)); -- 
    -- CP-element group 74:  branch  transition  place  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	70 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (13) 
      -- CP-element group 74: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540__exit__
      -- CP-element group 74: 	 branch_block_stmt_2214/if_stmt_2541__entry__
      -- CP-element group 74: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/$exit
      -- CP-element group 74: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2534_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2534_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2214/assign_stmt_2510_to_assign_stmt_2540/type_cast_2534_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_2214/if_stmt_2541_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2214/if_stmt_2541_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_2214/if_stmt_2541_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_2214/if_stmt_2541_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_2214/R_cmp122_2542_place
      -- CP-element group 74: 	 branch_block_stmt_2214/if_stmt_2541_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_2214/if_stmt_2541_else_link/$entry
      -- 
    ca_6404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2534_inst_ack_1, ack => convTransposeC_CP_5763_elements(74)); -- 
    branch_req_6412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(74), ack => if_stmt_2541_branch_req_0); -- 
    -- CP-element group 75:  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_2214/merge_stmt_2575__exit__
      -- CP-element group 75: 	 branch_block_stmt_2214/assign_stmt_2580__entry__
      -- CP-element group 75: 	 branch_block_stmt_2214/if_stmt_2541_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_2214/if_stmt_2541_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_2214/ifx_xelse_whilex_xend
      -- CP-element group 75: 	 branch_block_stmt_2214/assign_stmt_2580/$entry
      -- CP-element group 75: 	 branch_block_stmt_2214/assign_stmt_2580/WPIPE_Block2_done_2577_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_2214/assign_stmt_2580/WPIPE_Block2_done_2577_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_2214/assign_stmt_2580/WPIPE_Block2_done_2577_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_2214/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_2214/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_2214/merge_stmt_2575_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_2214/merge_stmt_2575_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_2214/merge_stmt_2575_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_2214/merge_stmt_2575_PhiAck/dummy
      -- 
    if_choice_transition_6417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2541_branch_ack_1, ack => convTransposeC_CP_5763_elements(75)); -- 
    req_6437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(75), ack => WPIPE_Block2_done_2577_inst_req_0); -- 
    -- CP-element group 76:  fork  transition  place  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	105 
    -- CP-element group 76: 	106 
    -- CP-element group 76: 	107 
    -- CP-element group 76: 	109 
    -- CP-element group 76: 	110 
    -- CP-element group 76:  members (22) 
      -- CP-element group 76: 	 branch_block_stmt_2214/if_stmt_2541_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_2214/if_stmt_2541_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2548/$entry
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/$entry
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/$entry
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/Update/cr
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2561/$entry
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2564/$entry
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2564/SplitProtocol/$entry
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2564/SplitProtocol/Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2564/SplitProtocol/Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2564/SplitProtocol/Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2564/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2541_branch_ack_0, ack => convTransposeC_CP_5763_elements(76)); -- 
    rr_6647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(76), ack => type_cast_2558_inst_req_0); -- 
    cr_6652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(76), ack => type_cast_2558_inst_req_1); -- 
    rr_6670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(76), ack => type_cast_2564_inst_req_0); -- 
    cr_6675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(76), ack => type_cast_2564_inst_req_1); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_2214/assign_stmt_2580/WPIPE_Block2_done_2577_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_2214/assign_stmt_2580/WPIPE_Block2_done_2577_update_start_
      -- CP-element group 77: 	 branch_block_stmt_2214/assign_stmt_2580/WPIPE_Block2_done_2577_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_2214/assign_stmt_2580/WPIPE_Block2_done_2577_Sample/ack
      -- CP-element group 77: 	 branch_block_stmt_2214/assign_stmt_2580/WPIPE_Block2_done_2577_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_2214/assign_stmt_2580/WPIPE_Block2_done_2577_Update/req
      -- 
    ack_6438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2577_inst_ack_0, ack => convTransposeC_CP_5763_elements(77)); -- 
    req_6442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(77), ack => WPIPE_Block2_done_2577_inst_req_1); -- 
    -- CP-element group 78:  transition  place  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (16) 
      -- CP-element group 78: 	 $exit
      -- CP-element group 78: 	 branch_block_stmt_2214/$exit
      -- CP-element group 78: 	 branch_block_stmt_2214/branch_block_stmt_2214__exit__
      -- CP-element group 78: 	 branch_block_stmt_2214/assign_stmt_2580__exit__
      -- CP-element group 78: 	 branch_block_stmt_2214/return__
      -- CP-element group 78: 	 branch_block_stmt_2214/merge_stmt_2582__exit__
      -- CP-element group 78: 	 branch_block_stmt_2214/assign_stmt_2580/$exit
      -- CP-element group 78: 	 branch_block_stmt_2214/assign_stmt_2580/WPIPE_Block2_done_2577_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_2214/assign_stmt_2580/WPIPE_Block2_done_2577_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_2214/assign_stmt_2580/WPIPE_Block2_done_2577_Update/ack
      -- CP-element group 78: 	 branch_block_stmt_2214/return___PhiReq/$entry
      -- CP-element group 78: 	 branch_block_stmt_2214/return___PhiReq/$exit
      -- CP-element group 78: 	 branch_block_stmt_2214/merge_stmt_2582_PhiReqMerge
      -- CP-element group 78: 	 branch_block_stmt_2214/merge_stmt_2582_PhiAck/$entry
      -- CP-element group 78: 	 branch_block_stmt_2214/merge_stmt_2582_PhiAck/$exit
      -- CP-element group 78: 	 branch_block_stmt_2214/merge_stmt_2582_PhiAck/dummy
      -- 
    ack_6443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2577_inst_ack_1, ack => convTransposeC_CP_5763_elements(78)); -- 
    -- CP-element group 79:  transition  output  delay-element  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	43 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	85 
    -- CP-element group 79:  members (4) 
      -- CP-element group 79: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2340/$exit
      -- CP-element group 79: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_sources/type_cast_2344_konst_delay_trans
      -- CP-element group 79: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_req
      -- 
    phi_stmt_2340_req_6454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2340_req_6454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(79), ack => phi_stmt_2340_req_0); -- 
    -- Element group convTransposeC_CP_5763_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convTransposeC_CP_5763_elements(43), ack => convTransposeC_CP_5763_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  transition  output  delay-element  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	43 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	85 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2347/$exit
      -- CP-element group 80: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_sources/type_cast_2353_konst_delay_trans
      -- CP-element group 80: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_req
      -- 
    phi_stmt_2347_req_6462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2347_req_6462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(80), ack => phi_stmt_2347_req_1); -- 
    -- Element group convTransposeC_CP_5763_elements(80) is a control-delay.
    cp_element_80_delay: control_delay_element  generic map(name => " 80_delay", delay_value => 1)  port map(req => convTransposeC_CP_5763_elements(43), ack => convTransposeC_CP_5763_elements(80), clk => clk, reset =>reset);
    -- CP-element group 81:  transition  output  delay-element  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	85 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2354/$exit
      -- CP-element group 81: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_sources/type_cast_2360_konst_delay_trans
      -- CP-element group 81: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_req
      -- 
    phi_stmt_2354_req_6470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2354_req_6470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(81), ack => phi_stmt_2354_req_1); -- 
    -- Element group convTransposeC_CP_5763_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convTransposeC_CP_5763_elements(43), ack => convTransposeC_CP_5763_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	43 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2366/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2366/SplitProtocol/Sample/ra
      -- 
    ra_6487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2366_inst_ack_0, ack => convTransposeC_CP_5763_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	43 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2366/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2366/SplitProtocol/Update/ca
      -- 
    ca_6492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2366_inst_ack_1, ack => convTransposeC_CP_5763_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2361/$exit
      -- CP-element group 84: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2366/$exit
      -- CP-element group 84: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2366/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_req
      -- 
    phi_stmt_2361_req_6493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2361_req_6493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(84), ack => phi_stmt_2361_req_1); -- 
    convTransposeC_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(82) & convTransposeC_CP_5763_elements(83);
      gj_convTransposeC_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	79 
    -- CP-element group 85: 	80 
    -- CP-element group 85: 	81 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	99 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2214/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(79) & convTransposeC_CP_5763_elements(80) & convTransposeC_CP_5763_elements(81) & convTransposeC_CP_5763_elements(84);
      gj_convTransposeC_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_sources/type_cast_2346/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_sources/type_cast_2346/SplitProtocol/Sample/ra
      -- 
    ra_6513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2346_inst_ack_0, ack => convTransposeC_CP_5763_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	1 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_sources/type_cast_2346/SplitProtocol/Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_sources/type_cast_2346/SplitProtocol/Update/ca
      -- 
    ca_6518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2346_inst_ack_1, ack => convTransposeC_CP_5763_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	98 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2340/$exit
      -- CP-element group 88: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_sources/$exit
      -- CP-element group 88: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_sources/type_cast_2346/$exit
      -- CP-element group 88: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_sources/type_cast_2346/SplitProtocol/$exit
      -- CP-element group 88: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2340/phi_stmt_2340_req
      -- 
    phi_stmt_2340_req_6519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2340_req_6519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(88), ack => phi_stmt_2340_req_1); -- 
    convTransposeC_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(86) & convTransposeC_CP_5763_elements(87);
      gj_convTransposeC_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_sources/type_cast_2350/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_sources/type_cast_2350/SplitProtocol/Sample/ra
      -- 
    ra_6536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2350_inst_ack_0, ack => convTransposeC_CP_5763_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	1 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_sources/type_cast_2350/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_sources/type_cast_2350/SplitProtocol/Update/ca
      -- 
    ca_6541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2350_inst_ack_1, ack => convTransposeC_CP_5763_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	98 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2347/$exit
      -- CP-element group 91: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_sources/type_cast_2350/$exit
      -- CP-element group 91: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_sources/type_cast_2350/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2347/phi_stmt_2347_req
      -- 
    phi_stmt_2347_req_6542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2347_req_6542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(91), ack => phi_stmt_2347_req_0); -- 
    convTransposeC_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(89) & convTransposeC_CP_5763_elements(90);
      gj_convTransposeC_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_sources/type_cast_2357/SplitProtocol/Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_sources/type_cast_2357/SplitProtocol/Sample/ra
      -- 
    ra_6559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2357_inst_ack_0, ack => convTransposeC_CP_5763_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	1 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_sources/type_cast_2357/SplitProtocol/Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_sources/type_cast_2357/SplitProtocol/Update/ca
      -- 
    ca_6564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2357_inst_ack_1, ack => convTransposeC_CP_5763_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	98 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2354/$exit
      -- CP-element group 94: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_sources/$exit
      -- CP-element group 94: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_sources/type_cast_2357/$exit
      -- CP-element group 94: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_sources/type_cast_2357/SplitProtocol/$exit
      -- CP-element group 94: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2354/phi_stmt_2354_req
      -- 
    phi_stmt_2354_req_6565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2354_req_6565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(94), ack => phi_stmt_2354_req_0); -- 
    convTransposeC_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(92) & convTransposeC_CP_5763_elements(93);
      gj_convTransposeC_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	1 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2364/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2364/SplitProtocol/Sample/ra
      -- 
    ra_6582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2364_inst_ack_0, ack => convTransposeC_CP_5763_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	1 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2364/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2364/SplitProtocol/Update/ca
      -- 
    ca_6587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2364_inst_ack_1, ack => convTransposeC_CP_5763_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2361/$exit
      -- CP-element group 97: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2364/$exit
      -- CP-element group 97: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_sources/type_cast_2364/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/phi_stmt_2361/phi_stmt_2361_req
      -- 
    phi_stmt_2361_req_6588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2361_req_6588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(97), ack => phi_stmt_2361_req_0); -- 
    convTransposeC_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(95) & convTransposeC_CP_5763_elements(96);
      gj_convTransposeC_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	88 
    -- CP-element group 98: 	91 
    -- CP-element group 98: 	94 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2214/ifx_xend133_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(88) & convTransposeC_CP_5763_elements(91) & convTransposeC_CP_5763_elements(94) & convTransposeC_CP_5763_elements(97);
      gj_convTransposeC_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  fork  transition  place  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	85 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	101 
    -- CP-element group 99: 	102 
    -- CP-element group 99: 	103 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2214/merge_stmt_2339_PhiReqMerge
      -- CP-element group 99: 	 branch_block_stmt_2214/merge_stmt_2339_PhiAck/$entry
      -- 
    convTransposeC_CP_5763_elements(99) <= OrReduce(convTransposeC_CP_5763_elements(85) & convTransposeC_CP_5763_elements(98));
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	104 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_2214/merge_stmt_2339_PhiAck/phi_stmt_2340_ack
      -- 
    phi_stmt_2340_ack_6593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2340_ack_0, ack => convTransposeC_CP_5763_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_2214/merge_stmt_2339_PhiAck/phi_stmt_2347_ack
      -- 
    phi_stmt_2347_ack_6594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2347_ack_0, ack => convTransposeC_CP_5763_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_2214/merge_stmt_2339_PhiAck/phi_stmt_2354_ack
      -- 
    phi_stmt_2354_ack_6595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2354_ack_0, ack => convTransposeC_CP_5763_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_2214/merge_stmt_2339_PhiAck/phi_stmt_2361_ack
      -- 
    phi_stmt_2361_ack_6596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2361_ack_0, ack => convTransposeC_CP_5763_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  place  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	100 
    -- CP-element group 104: 	101 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	44 
    -- CP-element group 104: 	45 
    -- CP-element group 104: 	46 
    -- CP-element group 104: 	47 
    -- CP-element group 104: 	48 
    -- CP-element group 104: 	49 
    -- CP-element group 104: 	50 
    -- CP-element group 104: 	51 
    -- CP-element group 104: 	53 
    -- CP-element group 104: 	55 
    -- CP-element group 104: 	57 
    -- CP-element group 104: 	60 
    -- CP-element group 104: 	62 
    -- CP-element group 104: 	65 
    -- CP-element group 104: 	66 
    -- CP-element group 104: 	67 
    -- CP-element group 104:  members (56) 
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2401_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2214/merge_stmt_2339__exit__
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489__entry__
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2401_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2401_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2401_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2401_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2401_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2405_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2405_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2405_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2405_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2405_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2405_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2409_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2409_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2409_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2409_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2409_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2409_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2439_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2439_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2439_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2439_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2439_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2439_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2446_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2445_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2446_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2446_complete/req
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2450_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2469_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_final_index_sum_regn_update_start
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_final_index_sum_regn_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/array_obj_ref_2468_final_index_sum_regn_Update/req
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2469_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/addr_of_2469_complete/req
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Update/word_access_complete/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Update/word_access_complete/word_0/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/ptr_deref_2472_Update/word_access_complete/word_0/cr
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2477_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2477_update_start_
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2477_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2477_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2477_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_2214/assign_stmt_2373_to_assign_stmt_2489/type_cast_2477_Update/cr
      -- CP-element group 104: 	 branch_block_stmt_2214/merge_stmt_2339_PhiAck/$exit
      -- 
    rr_6097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2401_inst_req_0); -- 
    cr_6102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2401_inst_req_1); -- 
    rr_6111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2405_inst_req_0); -- 
    cr_6116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2405_inst_req_1); -- 
    rr_6125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2409_inst_req_0); -- 
    cr_6130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2409_inst_req_1); -- 
    rr_6139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2439_inst_req_0); -- 
    cr_6144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2439_inst_req_1); -- 
    req_6175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => array_obj_ref_2445_index_offset_req_1); -- 
    req_6190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => addr_of_2446_final_reg_req_1); -- 
    cr_6235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => ptr_deref_2450_load_0_req_1); -- 
    req_6271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => array_obj_ref_2468_index_offset_req_1); -- 
    req_6286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => addr_of_2469_final_reg_req_1); -- 
    cr_6336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => ptr_deref_2472_store_0_req_1); -- 
    rr_6345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2477_inst_req_0); -- 
    cr_6350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(104), ack => type_cast_2477_inst_req_1); -- 
    convTransposeC_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(100) & convTransposeC_CP_5763_elements(101) & convTransposeC_CP_5763_elements(102) & convTransposeC_CP_5763_elements(103);
      gj_convTransposeC_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  output  delay-element  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	76 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	112 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2548/$exit
      -- CP-element group 105: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_sources/$exit
      -- CP-element group 105: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_sources/type_cast_2554_konst_delay_trans
      -- CP-element group 105: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_req
      -- 
    phi_stmt_2548_req_6631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2548_req_6631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(105), ack => phi_stmt_2548_req_1); -- 
    -- Element group convTransposeC_CP_5763_elements(105) is a control-delay.
    cp_element_105_delay: control_delay_element  generic map(name => " 105_delay", delay_value => 1)  port map(req => convTransposeC_CP_5763_elements(76), ack => convTransposeC_CP_5763_elements(105), clk => clk, reset =>reset);
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	76 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/Sample/ra
      -- 
    ra_6648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2558_inst_ack_0, ack => convTransposeC_CP_5763_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	76 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/Update/ca
      -- 
    ca_6653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2558_inst_ack_1, ack => convTransposeC_CP_5763_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/$exit
      -- CP-element group 108: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/$exit
      -- CP-element group 108: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2558/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_req
      -- 
    phi_stmt_2555_req_6654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2555_req_6654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(108), ack => phi_stmt_2555_req_0); -- 
    convTransposeC_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(106) & convTransposeC_CP_5763_elements(107);
      gj_convTransposeC_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	76 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2564/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2564/SplitProtocol/Sample/ra
      -- 
    ra_6671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2564_inst_ack_0, ack => convTransposeC_CP_5763_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	76 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2564/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2564/SplitProtocol/Update/ca
      -- 
    ca_6676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2564_inst_ack_1, ack => convTransposeC_CP_5763_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2561/$exit
      -- CP-element group 111: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2564/$exit
      -- CP-element group 111: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2564/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_req
      -- 
    phi_stmt_2561_req_6677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2561_req_6677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(111), ack => phi_stmt_2561_req_0); -- 
    convTransposeC_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(109) & convTransposeC_CP_5763_elements(110);
      gj_convTransposeC_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	105 
    -- CP-element group 112: 	108 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	123 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2214/ifx_xelse_ifx_xend133_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(105) & convTransposeC_CP_5763_elements(108) & convTransposeC_CP_5763_elements(111);
      gj_convTransposeC_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	69 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_sources/type_cast_2551/SplitProtocol/Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_sources/type_cast_2551/SplitProtocol/Sample/ra
      -- 
    ra_6697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2551_inst_ack_0, ack => convTransposeC_CP_5763_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	69 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_sources/type_cast_2551/SplitProtocol/Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_sources/type_cast_2551/SplitProtocol/Update/ca
      -- 
    ca_6702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2551_inst_ack_1, ack => convTransposeC_CP_5763_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	122 
    -- CP-element group 115:  members (5) 
      -- CP-element group 115: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2548/$exit
      -- CP-element group 115: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_sources/$exit
      -- CP-element group 115: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_sources/type_cast_2551/$exit
      -- CP-element group 115: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_sources/type_cast_2551/SplitProtocol/$exit
      -- CP-element group 115: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2548/phi_stmt_2548_req
      -- 
    phi_stmt_2548_req_6703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2548_req_6703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(115), ack => phi_stmt_2548_req_0); -- 
    convTransposeC_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(113) & convTransposeC_CP_5763_elements(114);
      gj_convTransposeC_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/Sample/ra
      -- 
    ra_6720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2560_inst_ack_0, ack => convTransposeC_CP_5763_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	69 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/Update/ca
      -- 
    ca_6725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2560_inst_ack_1, ack => convTransposeC_CP_5763_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	122 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/$exit
      -- CP-element group 118: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/$exit
      -- CP-element group 118: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/$exit
      -- CP-element group 118: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_sources/type_cast_2560/SplitProtocol/$exit
      -- CP-element group 118: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2555/phi_stmt_2555_req
      -- 
    phi_stmt_2555_req_6726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2555_req_6726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(118), ack => phi_stmt_2555_req_1); -- 
    convTransposeC_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(116) & convTransposeC_CP_5763_elements(117);
      gj_convTransposeC_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	69 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2566/SplitProtocol/Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2566/SplitProtocol/Sample/ra
      -- 
    ra_6743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2566_inst_ack_0, ack => convTransposeC_CP_5763_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	69 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2566/SplitProtocol/Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2566/SplitProtocol/Update/ca
      -- 
    ca_6748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2566_inst_ack_1, ack => convTransposeC_CP_5763_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (5) 
      -- CP-element group 121: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2561/$exit
      -- CP-element group 121: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/$exit
      -- CP-element group 121: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2566/$exit
      -- CP-element group 121: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_sources/type_cast_2566/SplitProtocol/$exit
      -- CP-element group 121: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/phi_stmt_2561/phi_stmt_2561_req
      -- 
    phi_stmt_2561_req_6749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2561_req_6749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5763_elements(121), ack => phi_stmt_2561_req_1); -- 
    convTransposeC_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(119) & convTransposeC_CP_5763_elements(120);
      gj_convTransposeC_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	115 
    -- CP-element group 122: 	118 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2214/ifx_xthen_ifx_xend133_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(115) & convTransposeC_CP_5763_elements(118) & convTransposeC_CP_5763_elements(121);
      gj_convTransposeC_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	112 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_2214/merge_stmt_2547_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_2214/merge_stmt_2547_PhiAck/$entry
      -- 
    convTransposeC_CP_5763_elements(123) <= OrReduce(convTransposeC_CP_5763_elements(112) & convTransposeC_CP_5763_elements(122));
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	127 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_2214/merge_stmt_2547_PhiAck/phi_stmt_2548_ack
      -- 
    phi_stmt_2548_ack_6754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2548_ack_0, ack => convTransposeC_CP_5763_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_2214/merge_stmt_2547_PhiAck/phi_stmt_2555_ack
      -- 
    phi_stmt_2555_ack_6755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2555_ack_0, ack => convTransposeC_CP_5763_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_2214/merge_stmt_2547_PhiAck/phi_stmt_2561_ack
      -- 
    phi_stmt_2561_ack_6756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2561_ack_0, ack => convTransposeC_CP_5763_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	124 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_2214/merge_stmt_2547_PhiAck/$exit
      -- 
    convTransposeC_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5763_elements(124) & convTransposeC_CP_5763_elements(125) & convTransposeC_CP_5763_elements(126);
      gj_convTransposeC_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5763_elements(127), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom86_2467_resized : std_logic_vector(13 downto 0);
    signal R_idxprom86_2467_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2444_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2444_scaled : std_logic_vector(13 downto 0);
    signal add121_2337 : std_logic_vector(31 downto 0);
    signal add45_2288 : std_logic_vector(15 downto 0);
    signal add58_2299 : std_logic_vector(15 downto 0);
    signal add77_2420 : std_logic_vector(63 downto 0);
    signal add79_2430 : std_logic_vector(63 downto 0);
    signal add91_2484 : std_logic_vector(31 downto 0);
    signal add98_2502 : std_logic_vector(15 downto 0);
    signal add_2266 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2378 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2445_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2445_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2445_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2445_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2445_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2445_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2468_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2468_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2468_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2468_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2468_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2468_root_address : std_logic_vector(13 downto 0);
    signal arrayidx82_2447 : std_logic_vector(31 downto 0);
    signal arrayidx87_2470 : std_logic_vector(31 downto 0);
    signal call11_2235 : std_logic_vector(15 downto 0);
    signal call13_2238 : std_logic_vector(15 downto 0);
    signal call14_2241 : std_logic_vector(15 downto 0);
    signal call15_2244 : std_logic_vector(15 downto 0);
    signal call16_2257 : std_logic_vector(15 downto 0);
    signal call18_2269 : std_logic_vector(15 downto 0);
    signal call1_2220 : std_logic_vector(15 downto 0);
    signal call20_2272 : std_logic_vector(15 downto 0);
    signal call22_2275 : std_logic_vector(15 downto 0);
    signal call3_2223 : std_logic_vector(15 downto 0);
    signal call5_2226 : std_logic_vector(15 downto 0);
    signal call7_2229 : std_logic_vector(15 downto 0);
    signal call9_2232 : std_logic_vector(15 downto 0);
    signal call_2217 : std_logic_vector(15 downto 0);
    signal cmp106_2515 : std_logic_vector(0 downto 0);
    signal cmp122_2540 : std_logic_vector(0 downto 0);
    signal cmp_2489 : std_logic_vector(0 downto 0);
    signal conv112_2535 : std_logic_vector(31 downto 0);
    signal conv115_2320 : std_logic_vector(31 downto 0);
    signal conv17_2261 : std_logic_vector(31 downto 0);
    signal conv65_2402 : std_logic_vector(63 downto 0);
    signal conv68_2308 : std_logic_vector(63 downto 0);
    signal conv70_2406 : std_logic_vector(63 downto 0);
    signal conv73_2312 : std_logic_vector(63 downto 0);
    signal conv75_2410 : std_logic_vector(63 downto 0);
    signal conv90_2478 : std_logic_vector(31 downto 0);
    signal conv94_2316 : std_logic_vector(31 downto 0);
    signal conv_2248 : std_logic_vector(31 downto 0);
    signal idxprom86_2463 : std_logic_vector(63 downto 0);
    signal idxprom_2440 : std_logic_vector(63 downto 0);
    signal inc110_2519 : std_logic_vector(15 downto 0);
    signal inc110x_xinput_dim0x_x2_2524 : std_logic_vector(15 downto 0);
    signal inc_2510 : std_logic_vector(15 downto 0);
    signal indvar_2340 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2573 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2561 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2361 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2555 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2354 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2531 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2548 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2347 : std_logic_vector(15 downto 0);
    signal mul54_2393 : std_logic_vector(15 downto 0);
    signal mul76_2415 : std_logic_vector(63 downto 0);
    signal mul78_2425 : std_logic_vector(63 downto 0);
    signal mul_2383 : std_logic_vector(15 downto 0);
    signal ptr_deref_2450_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2450_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2450_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2450_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2450_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2472_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2472_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2472_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2472_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2472_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2472_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2254 : std_logic_vector(31 downto 0);
    signal shr116137_2326 : std_logic_vector(31 downto 0);
    signal shr120138_2332 : std_logic_vector(31 downto 0);
    signal shr136_2282 : std_logic_vector(15 downto 0);
    signal shr81_2436 : std_logic_vector(31 downto 0);
    signal shr85_2457 : std_logic_vector(63 downto 0);
    signal sub48_2388 : std_logic_vector(15 downto 0);
    signal sub61_2304 : std_logic_vector(15 downto 0);
    signal sub62_2398 : std_logic_vector(15 downto 0);
    signal sub_2293 : std_logic_vector(15 downto 0);
    signal tmp1_2373 : std_logic_vector(31 downto 0);
    signal tmp83_2451 : std_logic_vector(63 downto 0);
    signal type_cast_2252_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2280_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2286_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2297_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2324_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2330_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2344_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2346_wire : std_logic_vector(31 downto 0);
    signal type_cast_2350_wire : std_logic_vector(15 downto 0);
    signal type_cast_2353_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2357_wire : std_logic_vector(15 downto 0);
    signal type_cast_2360_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2364_wire : std_logic_vector(15 downto 0);
    signal type_cast_2366_wire : std_logic_vector(15 downto 0);
    signal type_cast_2371_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2434_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2455_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2461_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2482_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2500_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2508_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2528_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2551_wire : std_logic_vector(15 downto 0);
    signal type_cast_2554_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2558_wire : std_logic_vector(15 downto 0);
    signal type_cast_2560_wire : std_logic_vector(15 downto 0);
    signal type_cast_2564_wire : std_logic_vector(15 downto 0);
    signal type_cast_2566_wire : std_logic_vector(15 downto 0);
    signal type_cast_2571_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2579_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2445_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2445_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2445_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2445_resized_base_address <= "00000000000000";
    array_obj_ref_2468_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2468_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2468_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2468_resized_base_address <= "00000000000000";
    ptr_deref_2450_word_offset_0 <= "00000000000000";
    ptr_deref_2472_word_offset_0 <= "00000000000000";
    type_cast_2252_wire_constant <= "00000000000000000000000000010000";
    type_cast_2280_wire_constant <= "0000000000000001";
    type_cast_2286_wire_constant <= "1111111111111111";
    type_cast_2297_wire_constant <= "1111111111111111";
    type_cast_2324_wire_constant <= "00000000000000000000000000000010";
    type_cast_2330_wire_constant <= "00000000000000000000000000000001";
    type_cast_2344_wire_constant <= "00000000000000000000000000000000";
    type_cast_2353_wire_constant <= "0000000000000000";
    type_cast_2360_wire_constant <= "0000000000000000";
    type_cast_2371_wire_constant <= "00000000000000000000000000000100";
    type_cast_2434_wire_constant <= "00000000000000000000000000000010";
    type_cast_2455_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2461_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2482_wire_constant <= "00000000000000000000000000000100";
    type_cast_2500_wire_constant <= "0000000000000100";
    type_cast_2508_wire_constant <= "0000000000000001";
    type_cast_2528_wire_constant <= "0000000000000000";
    type_cast_2554_wire_constant <= "0000000000000000";
    type_cast_2571_wire_constant <= "00000000000000000000000000000001";
    type_cast_2579_wire_constant <= "0000000000000001";
    phi_stmt_2340: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2344_wire_constant & type_cast_2346_wire;
      req <= phi_stmt_2340_req_0 & phi_stmt_2340_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2340",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2340_ack_0,
          idata => idata,
          odata => indvar_2340,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2340
    phi_stmt_2347: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2350_wire & type_cast_2353_wire_constant;
      req <= phi_stmt_2347_req_0 & phi_stmt_2347_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2347",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2347_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2347,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2347
    phi_stmt_2354: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2357_wire & type_cast_2360_wire_constant;
      req <= phi_stmt_2354_req_0 & phi_stmt_2354_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2354",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2354_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2354,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2354
    phi_stmt_2361: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2364_wire & type_cast_2366_wire;
      req <= phi_stmt_2361_req_0 & phi_stmt_2361_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2361",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2361_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2361,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2361
    phi_stmt_2548: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2551_wire & type_cast_2554_wire_constant;
      req <= phi_stmt_2548_req_0 & phi_stmt_2548_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2548",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2548_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2548,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2548
    phi_stmt_2555: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2558_wire & type_cast_2560_wire;
      req <= phi_stmt_2555_req_0 & phi_stmt_2555_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2555",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2555_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2555,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2555
    phi_stmt_2561: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2564_wire & type_cast_2566_wire;
      req <= phi_stmt_2561_req_0 & phi_stmt_2561_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2561",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2561_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2561,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2561
    -- flow-through select operator MUX_2530_inst
    input_dim1x_x2_2531 <= type_cast_2528_wire_constant when (cmp106_2515(0) /=  '0') else inc_2510;
    addr_of_2446_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2446_final_reg_req_0;
      addr_of_2446_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2446_final_reg_req_1;
      addr_of_2446_final_reg_ack_1<= rack(0);
      addr_of_2446_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2446_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2445_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx82_2447,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2469_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2469_final_reg_req_0;
      addr_of_2469_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2469_final_reg_req_1;
      addr_of_2469_final_reg_ack_1<= rack(0);
      addr_of_2469_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2469_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2468_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2470,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2247_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2247_inst_req_0;
      type_cast_2247_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2247_inst_req_1;
      type_cast_2247_inst_ack_1<= rack(0);
      type_cast_2247_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2247_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2244,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2248,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2260_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2260_inst_req_0;
      type_cast_2260_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2260_inst_req_1;
      type_cast_2260_inst_ack_1<= rack(0);
      type_cast_2260_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2260_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2257,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2261,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2307_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2307_inst_req_0;
      type_cast_2307_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2307_inst_req_1;
      type_cast_2307_inst_ack_1<= rack(0);
      type_cast_2307_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2307_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2275,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_2308,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2311_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2311_inst_req_0;
      type_cast_2311_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2311_inst_req_1;
      type_cast_2311_inst_ack_1<= rack(0);
      type_cast_2311_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2311_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2272,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2312,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2315_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2315_inst_req_0;
      type_cast_2315_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2315_inst_req_1;
      type_cast_2315_inst_ack_1<= rack(0);
      type_cast_2315_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2315_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2223,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv94_2316,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2319_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2319_inst_req_0;
      type_cast_2319_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2319_inst_req_1;
      type_cast_2319_inst_ack_1<= rack(0);
      type_cast_2319_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2319_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_2217,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_2320,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2346_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2346_inst_req_0;
      type_cast_2346_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2346_inst_req_1;
      type_cast_2346_inst_ack_1<= rack(0);
      type_cast_2346_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2346_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2573,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2346_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2350_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2350_inst_req_0;
      type_cast_2350_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2350_inst_req_1;
      type_cast_2350_inst_ack_1<= rack(0);
      type_cast_2350_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2350_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2548,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2350_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2357_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2357_inst_req_0;
      type_cast_2357_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2357_inst_req_1;
      type_cast_2357_inst_ack_1<= rack(0);
      type_cast_2357_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2357_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2555,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2357_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2364_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2364_inst_req_0;
      type_cast_2364_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2364_inst_req_1;
      type_cast_2364_inst_ack_1<= rack(0);
      type_cast_2364_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2364_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2561,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2364_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2366_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2366_inst_req_0;
      type_cast_2366_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2366_inst_req_1;
      type_cast_2366_inst_ack_1<= rack(0);
      type_cast_2366_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2366_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr136_2282,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2366_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2401_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2401_inst_req_0;
      type_cast_2401_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2401_inst_req_1;
      type_cast_2401_inst_ack_1<= rack(0);
      type_cast_2401_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2401_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2347,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2402,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2405_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2405_inst_req_0;
      type_cast_2405_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2405_inst_req_1;
      type_cast_2405_inst_ack_1<= rack(0);
      type_cast_2405_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2405_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub62_2398,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2406,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2409_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2409_inst_req_0;
      type_cast_2409_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2409_inst_req_1;
      type_cast_2409_inst_ack_1<= rack(0);
      type_cast_2409_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2409_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub48_2388,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2410,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2439_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2439_inst_req_0;
      type_cast_2439_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2439_inst_req_1;
      type_cast_2439_inst_ack_1<= rack(0);
      type_cast_2439_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2439_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr81_2436,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2440,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2477_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2477_inst_req_0;
      type_cast_2477_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2477_inst_req_1;
      type_cast_2477_inst_ack_1<= rack(0);
      type_cast_2477_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2477_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2347,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_2478,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2518_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2518_inst_req_0;
      type_cast_2518_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2518_inst_req_1;
      type_cast_2518_inst_ack_1<= rack(0);
      type_cast_2518_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2518_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp106_2515,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc110_2519,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2534_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2534_inst_req_0;
      type_cast_2534_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2534_inst_req_1;
      type_cast_2534_inst_ack_1<= rack(0);
      type_cast_2534_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2534_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2524,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv112_2535,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2551_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2551_inst_req_0;
      type_cast_2551_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2551_inst_req_1;
      type_cast_2551_inst_ack_1<= rack(0);
      type_cast_2551_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2551_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add98_2502,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2551_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2558_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2558_inst_req_0;
      type_cast_2558_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2558_inst_req_1;
      type_cast_2558_inst_ack_1<= rack(0);
      type_cast_2558_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2558_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2531,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2558_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2560_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2560_inst_req_0;
      type_cast_2560_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2560_inst_req_1;
      type_cast_2560_inst_ack_1<= rack(0);
      type_cast_2560_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2560_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2354,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2560_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2564_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2564_inst_req_0;
      type_cast_2564_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2564_inst_req_1;
      type_cast_2564_inst_ack_1<= rack(0);
      type_cast_2564_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2564_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc110x_xinput_dim0x_x2_2524,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2564_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2566_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2566_inst_req_0;
      type_cast_2566_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2566_inst_req_1;
      type_cast_2566_inst_ack_1<= rack(0);
      type_cast_2566_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2566_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2361,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2566_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2445_index_1_rename
    process(R_idxprom_2444_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2444_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2444_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2445_index_1_resize
    process(idxprom_2440) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2440;
      ov := iv(13 downto 0);
      R_idxprom_2444_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2445_root_address_inst
    process(array_obj_ref_2445_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2445_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2445_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2468_index_1_rename
    process(R_idxprom86_2467_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom86_2467_resized;
      ov(13 downto 0) := iv;
      R_idxprom86_2467_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2468_index_1_resize
    process(idxprom86_2463) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom86_2463;
      ov := iv(13 downto 0);
      R_idxprom86_2467_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2468_root_address_inst
    process(array_obj_ref_2468_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2468_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2468_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2450_addr_0
    process(ptr_deref_2450_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2450_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2450_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2450_base_resize
    process(arrayidx82_2447) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx82_2447;
      ov := iv(13 downto 0);
      ptr_deref_2450_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2450_gather_scatter
    process(ptr_deref_2450_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2450_data_0;
      ov(63 downto 0) := iv;
      tmp83_2451 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2450_root_address_inst
    process(ptr_deref_2450_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2450_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2450_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2472_addr_0
    process(ptr_deref_2472_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2472_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2472_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2472_base_resize
    process(arrayidx87_2470) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2470;
      ov := iv(13 downto 0);
      ptr_deref_2472_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2472_gather_scatter
    process(tmp83_2451) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp83_2451;
      ov(63 downto 0) := iv;
      ptr_deref_2472_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2472_root_address_inst
    process(ptr_deref_2472_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2472_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2472_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2490_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2489;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2490_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2490_branch_req_0,
          ack0 => if_stmt_2490_branch_ack_0,
          ack1 => if_stmt_2490_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2541_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp122_2540;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2541_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2541_branch_req_0,
          ack0 => if_stmt_2541_branch_ack_0,
          ack1 => if_stmt_2541_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2287_inst
    process(call7_2229) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2229, type_cast_2286_wire_constant, tmp_var);
      add45_2288 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2298_inst
    process(call9_2232) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2232, type_cast_2297_wire_constant, tmp_var);
      add58_2299 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2387_inst
    process(sub_2293, mul_2383) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2293, mul_2383, tmp_var);
      sub48_2388 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2397_inst
    process(sub61_2304, mul54_2393) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub61_2304, mul54_2393, tmp_var);
      sub62_2398 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2501_inst
    process(input_dim2x_x1_2347) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2347, type_cast_2500_wire_constant, tmp_var);
      add98_2502 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2509_inst
    process(input_dim1x_x1_2354) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2354, type_cast_2508_wire_constant, tmp_var);
      inc_2510 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2523_inst
    process(inc110_2519, input_dim0x_x2_2361) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc110_2519, input_dim0x_x2_2361, tmp_var);
      inc110x_xinput_dim0x_x2_2524 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2336_inst
    process(shr116137_2326, shr120138_2332) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr116137_2326, shr120138_2332, tmp_var);
      add121_2337 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2377_inst
    process(add_2266, tmp1_2373) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2266, tmp1_2373, tmp_var);
      add_src_0x_x0_2378 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2483_inst
    process(conv90_2478) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv90_2478, type_cast_2482_wire_constant, tmp_var);
      add91_2484 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2572_inst
    process(indvar_2340) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2340, type_cast_2571_wire_constant, tmp_var);
      indvarx_xnext_2573 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2419_inst
    process(mul76_2415, conv70_2406) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul76_2415, conv70_2406, tmp_var);
      add77_2420 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2429_inst
    process(mul78_2425, conv65_2402) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul78_2425, conv65_2402, tmp_var);
      add79_2430 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2462_inst
    process(shr85_2457) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr85_2457, type_cast_2461_wire_constant, tmp_var);
      idxprom86_2463 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2514_inst
    process(inc_2510, call1_2220) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2510, call1_2220, tmp_var);
      cmp106_2515 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2539_inst
    process(conv112_2535, add121_2337) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv112_2535, add121_2337, tmp_var);
      cmp122_2540 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2281_inst
    process(call_2217) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2217, type_cast_2280_wire_constant, tmp_var);
      shr136_2282 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2325_inst
    process(conv115_2320) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_2320, type_cast_2324_wire_constant, tmp_var);
      shr116137_2326 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2331_inst
    process(conv115_2320) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv115_2320, type_cast_2330_wire_constant, tmp_var);
      shr120138_2332 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2435_inst
    process(add_src_0x_x0_2378) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2378, type_cast_2434_wire_constant, tmp_var);
      shr81_2436 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2456_inst
    process(add79_2430) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add79_2430, type_cast_2455_wire_constant, tmp_var);
      shr85_2457 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2382_inst
    process(input_dim0x_x2_2361, call13_2238) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2361, call13_2238, tmp_var);
      mul_2383 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2392_inst
    process(input_dim1x_x1_2354, call13_2238) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2354, call13_2238, tmp_var);
      mul54_2393 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2372_inst
    process(indvar_2340) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2340, type_cast_2371_wire_constant, tmp_var);
      tmp1_2373 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2414_inst
    process(conv75_2410, conv73_2312) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv75_2410, conv73_2312, tmp_var);
      mul76_2415 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2424_inst
    process(add77_2420, conv68_2308) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add77_2420, conv68_2308, tmp_var);
      mul78_2425 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2265_inst
    process(shl_2254, conv17_2261) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2254, conv17_2261, tmp_var);
      add_2266 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2253_inst
    process(conv_2248) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2248, type_cast_2252_wire_constant, tmp_var);
      shl_2254 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2292_inst
    process(add45_2288, call14_2241) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add45_2288, call14_2241, tmp_var);
      sub_2293 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2303_inst
    process(add58_2299, call14_2241) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add58_2299, call14_2241, tmp_var);
      sub61_2304 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2488_inst
    process(add91_2484, conv94_2316) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add91_2484, conv94_2316, tmp_var);
      cmp_2489 <= tmp_var; --
    end process;
    -- shared split operator group (31) : array_obj_ref_2445_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2444_scaled;
      array_obj_ref_2445_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2445_index_offset_req_0;
      array_obj_ref_2445_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2445_index_offset_req_1;
      array_obj_ref_2445_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : array_obj_ref_2468_index_offset 
    ApIntAdd_group_32: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom86_2467_scaled;
      array_obj_ref_2468_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2468_index_offset_req_0;
      array_obj_ref_2468_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2468_index_offset_req_1;
      array_obj_ref_2468_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_32_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared load operator group (0) : ptr_deref_2450_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2450_load_0_req_0;
      ptr_deref_2450_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2450_load_0_req_1;
      ptr_deref_2450_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2450_word_address_0;
      ptr_deref_2450_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2472_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2472_store_0_req_0;
      ptr_deref_2472_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2472_store_0_req_1;
      ptr_deref_2472_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2472_word_address_0;
      data_in <= ptr_deref_2472_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2268_inst RPIPE_Block2_start_2271_inst RPIPE_Block2_start_2256_inst RPIPE_Block2_start_2243_inst RPIPE_Block2_start_2240_inst RPIPE_Block2_start_2237_inst RPIPE_Block2_start_2234_inst RPIPE_Block2_start_2231_inst RPIPE_Block2_start_2228_inst RPIPE_Block2_start_2225_inst RPIPE_Block2_start_2222_inst RPIPE_Block2_start_2219_inst RPIPE_Block2_start_2274_inst RPIPE_Block2_start_2216_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block2_start_2268_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block2_start_2271_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block2_start_2256_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block2_start_2243_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block2_start_2240_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block2_start_2237_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block2_start_2234_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block2_start_2231_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block2_start_2228_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block2_start_2225_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block2_start_2222_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block2_start_2219_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block2_start_2274_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block2_start_2216_inst_req_0;
      RPIPE_Block2_start_2268_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block2_start_2271_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block2_start_2256_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block2_start_2243_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block2_start_2240_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block2_start_2237_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block2_start_2234_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block2_start_2231_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block2_start_2228_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block2_start_2225_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block2_start_2222_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block2_start_2219_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block2_start_2274_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block2_start_2216_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block2_start_2268_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block2_start_2271_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block2_start_2256_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block2_start_2243_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block2_start_2240_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block2_start_2237_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block2_start_2234_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block2_start_2231_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block2_start_2228_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block2_start_2225_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block2_start_2222_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block2_start_2219_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block2_start_2274_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block2_start_2216_inst_req_1;
      RPIPE_Block2_start_2268_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block2_start_2271_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block2_start_2256_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block2_start_2243_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block2_start_2240_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block2_start_2237_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block2_start_2234_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block2_start_2231_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block2_start_2228_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block2_start_2225_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block2_start_2222_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block2_start_2219_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block2_start_2274_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block2_start_2216_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call18_2269 <= data_out(223 downto 208);
      call20_2272 <= data_out(207 downto 192);
      call16_2257 <= data_out(191 downto 176);
      call15_2244 <= data_out(175 downto 160);
      call14_2241 <= data_out(159 downto 144);
      call13_2238 <= data_out(143 downto 128);
      call11_2235 <= data_out(127 downto 112);
      call9_2232 <= data_out(111 downto 96);
      call7_2229 <= data_out(95 downto 80);
      call5_2226 <= data_out(79 downto 64);
      call3_2223 <= data_out(63 downto 48);
      call1_2220 <= data_out(47 downto 32);
      call22_2275 <= data_out(31 downto 16);
      call_2217 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2577_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2577_inst_req_0;
      WPIPE_Block2_done_2577_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2577_inst_req_1;
      WPIPE_Block2_done_2577_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2579_wire_constant;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_6773_start: Boolean;
  signal convTransposeD_CP_6773_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block3_start_2646_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2646_inst_req_0 : boolean;
  signal type_cast_2632_inst_ack_0 : boolean;
  signal type_cast_2632_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2640_inst_req_0 : boolean;
  signal type_cast_2698_inst_ack_0 : boolean;
  signal addr_of_2808_final_reg_ack_1 : boolean;
  signal RPIPE_Block3_start_2646_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2646_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2640_inst_ack_1 : boolean;
  signal type_cast_2801_inst_req_1 : boolean;
  signal addr_of_2808_final_reg_req_1 : boolean;
  signal addr_of_2808_final_reg_req_0 : boolean;
  signal addr_of_2808_final_reg_ack_0 : boolean;
  signal RPIPE_Block3_start_2643_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2640_inst_ack_0 : boolean;
  signal type_cast_2771_inst_ack_1 : boolean;
  signal type_cast_2801_inst_req_0 : boolean;
  signal type_cast_2763_inst_req_0 : boolean;
  signal type_cast_2632_inst_ack_1 : boolean;
  signal type_cast_2763_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2643_inst_ack_1 : boolean;
  signal type_cast_2698_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2628_inst_req_0 : boolean;
  signal type_cast_2767_inst_req_1 : boolean;
  signal type_cast_2801_inst_ack_0 : boolean;
  signal type_cast_2690_inst_req_0 : boolean;
  signal type_cast_2619_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2628_inst_ack_0 : boolean;
  signal type_cast_2801_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2643_inst_ack_0 : boolean;
  signal type_cast_2767_inst_ack_1 : boolean;
  signal type_cast_2690_inst_ack_0 : boolean;
  signal type_cast_2694_inst_req_1 : boolean;
  signal type_cast_2698_inst_req_0 : boolean;
  signal type_cast_2767_inst_req_0 : boolean;
  signal type_cast_2694_inst_req_0 : boolean;
  signal type_cast_2771_inst_req_0 : boolean;
  signal type_cast_2690_inst_ack_1 : boolean;
  signal type_cast_2694_inst_ack_0 : boolean;
  signal type_cast_2694_inst_ack_1 : boolean;
  signal type_cast_2771_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2628_inst_req_1 : boolean;
  signal type_cast_2632_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2628_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2643_inst_req_1 : boolean;
  signal type_cast_2619_inst_req_1 : boolean;
  signal array_obj_ref_2807_index_offset_req_0 : boolean;
  signal type_cast_2767_inst_ack_0 : boolean;
  signal type_cast_2698_inst_ack_1 : boolean;
  signal array_obj_ref_2807_index_offset_ack_0 : boolean;
  signal array_obj_ref_2807_index_offset_req_1 : boolean;
  signal RPIPE_Block3_start_2640_inst_req_1 : boolean;
  signal type_cast_2771_inst_ack_0 : boolean;
  signal array_obj_ref_2807_index_offset_ack_1 : boolean;
  signal type_cast_2763_inst_req_1 : boolean;
  signal type_cast_2763_inst_ack_1 : boolean;
  signal type_cast_2690_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2588_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2588_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2588_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2588_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2591_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2591_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2591_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2591_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2594_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2594_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2594_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2594_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2597_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2597_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2597_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2597_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2600_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2600_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2600_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2600_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2603_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2603_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2603_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2603_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2606_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2606_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2606_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2606_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2609_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2609_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2609_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2609_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2612_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2612_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2612_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2612_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2615_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2615_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2615_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2615_inst_ack_1 : boolean;
  signal type_cast_2619_inst_req_0 : boolean;
  signal type_cast_2619_inst_ack_0 : boolean;
  signal ptr_deref_2812_load_0_req_0 : boolean;
  signal ptr_deref_2812_load_0_ack_0 : boolean;
  signal ptr_deref_2812_load_0_req_1 : boolean;
  signal ptr_deref_2812_load_0_ack_1 : boolean;
  signal array_obj_ref_2830_index_offset_req_0 : boolean;
  signal array_obj_ref_2830_index_offset_ack_0 : boolean;
  signal array_obj_ref_2830_index_offset_req_1 : boolean;
  signal array_obj_ref_2830_index_offset_ack_1 : boolean;
  signal addr_of_2831_final_reg_req_0 : boolean;
  signal addr_of_2831_final_reg_ack_0 : boolean;
  signal addr_of_2831_final_reg_req_1 : boolean;
  signal addr_of_2831_final_reg_ack_1 : boolean;
  signal ptr_deref_2834_store_0_req_0 : boolean;
  signal ptr_deref_2834_store_0_ack_0 : boolean;
  signal ptr_deref_2834_store_0_req_1 : boolean;
  signal ptr_deref_2834_store_0_ack_1 : boolean;
  signal type_cast_2839_inst_req_0 : boolean;
  signal type_cast_2839_inst_ack_0 : boolean;
  signal type_cast_2839_inst_req_1 : boolean;
  signal type_cast_2839_inst_ack_1 : boolean;
  signal if_stmt_2852_branch_req_0 : boolean;
  signal if_stmt_2852_branch_ack_1 : boolean;
  signal if_stmt_2852_branch_ack_0 : boolean;
  signal type_cast_2880_inst_req_0 : boolean;
  signal type_cast_2880_inst_ack_0 : boolean;
  signal type_cast_2880_inst_req_1 : boolean;
  signal type_cast_2880_inst_ack_1 : boolean;
  signal if_stmt_2899_branch_req_0 : boolean;
  signal if_stmt_2899_branch_ack_1 : boolean;
  signal if_stmt_2899_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_2935_inst_req_0 : boolean;
  signal WPIPE_Block3_done_2935_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_2935_inst_req_1 : boolean;
  signal WPIPE_Block3_done_2935_inst_ack_1 : boolean;
  signal phi_stmt_2702_req_0 : boolean;
  signal phi_stmt_2709_req_0 : boolean;
  signal phi_stmt_2716_req_0 : boolean;
  signal type_cast_2726_inst_req_0 : boolean;
  signal type_cast_2726_inst_ack_0 : boolean;
  signal type_cast_2726_inst_req_1 : boolean;
  signal type_cast_2726_inst_ack_1 : boolean;
  signal phi_stmt_2723_req_0 : boolean;
  signal type_cast_2708_inst_req_0 : boolean;
  signal type_cast_2708_inst_ack_0 : boolean;
  signal type_cast_2708_inst_req_1 : boolean;
  signal type_cast_2708_inst_ack_1 : boolean;
  signal phi_stmt_2702_req_1 : boolean;
  signal type_cast_2715_inst_req_0 : boolean;
  signal type_cast_2715_inst_ack_0 : boolean;
  signal type_cast_2715_inst_req_1 : boolean;
  signal type_cast_2715_inst_ack_1 : boolean;
  signal phi_stmt_2709_req_1 : boolean;
  signal type_cast_2722_inst_req_0 : boolean;
  signal type_cast_2722_inst_ack_0 : boolean;
  signal type_cast_2722_inst_req_1 : boolean;
  signal type_cast_2722_inst_ack_1 : boolean;
  signal phi_stmt_2716_req_1 : boolean;
  signal type_cast_2728_inst_req_0 : boolean;
  signal type_cast_2728_inst_ack_0 : boolean;
  signal type_cast_2728_inst_req_1 : boolean;
  signal type_cast_2728_inst_ack_1 : boolean;
  signal phi_stmt_2723_req_1 : boolean;
  signal phi_stmt_2702_ack_0 : boolean;
  signal phi_stmt_2709_ack_0 : boolean;
  signal phi_stmt_2716_ack_0 : boolean;
  signal phi_stmt_2723_ack_0 : boolean;
  signal phi_stmt_2906_req_1 : boolean;
  signal type_cast_2918_inst_req_0 : boolean;
  signal type_cast_2918_inst_ack_0 : boolean;
  signal type_cast_2918_inst_req_1 : boolean;
  signal type_cast_2918_inst_ack_1 : boolean;
  signal phi_stmt_2913_req_1 : boolean;
  signal type_cast_2924_inst_req_0 : boolean;
  signal type_cast_2924_inst_ack_0 : boolean;
  signal type_cast_2924_inst_req_1 : boolean;
  signal type_cast_2924_inst_ack_1 : boolean;
  signal phi_stmt_2919_req_1 : boolean;
  signal type_cast_2909_inst_req_0 : boolean;
  signal type_cast_2909_inst_ack_0 : boolean;
  signal type_cast_2909_inst_req_1 : boolean;
  signal type_cast_2909_inst_ack_1 : boolean;
  signal phi_stmt_2906_req_0 : boolean;
  signal type_cast_2916_inst_req_0 : boolean;
  signal type_cast_2916_inst_ack_0 : boolean;
  signal type_cast_2916_inst_req_1 : boolean;
  signal type_cast_2916_inst_ack_1 : boolean;
  signal phi_stmt_2913_req_0 : boolean;
  signal type_cast_2922_inst_req_0 : boolean;
  signal type_cast_2922_inst_ack_0 : boolean;
  signal type_cast_2922_inst_req_1 : boolean;
  signal type_cast_2922_inst_ack_1 : boolean;
  signal phi_stmt_2919_req_0 : boolean;
  signal phi_stmt_2906_ack_0 : boolean;
  signal phi_stmt_2913_ack_0 : boolean;
  signal phi_stmt_2919_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_6773_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6773_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_6773_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6773_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_6773: Block -- control-path 
    signal convTransposeD_CP_6773_elements: BooleanArray(123 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_6773_elements(0) <= convTransposeD_CP_6773_start;
    convTransposeD_CP_6773_symbol <= convTransposeD_CP_6773_elements(74);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	23 
    -- CP-element group 0: 	27 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2632_update_start_
      -- CP-element group 0: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2632_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2619_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2632_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2619_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2586/$entry
      -- CP-element group 0: 	 branch_block_stmt_2586/branch_block_stmt_2586__entry__
      -- CP-element group 0: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647__entry__
      -- CP-element group 0: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/$entry
      -- CP-element group 0: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2588_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2588_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2588_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2619_update_start_
      -- 
    cr_6994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(0), ack => type_cast_2632_inst_req_1); -- 
    cr_6966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(0), ack => type_cast_2619_inst_req_1); -- 
    rr_6821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(0), ack => RPIPE_Block3_start_2588_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	123 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	82 
    -- CP-element group 1: 	83 
    -- CP-element group 1: 	85 
    -- CP-element group 1: 	86 
    -- CP-element group 1: 	88 
    -- CP-element group 1: 	89 
    -- CP-element group 1: 	91 
    -- CP-element group 1: 	92 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2586/merge_stmt_2905__exit__
      -- CP-element group 1: 	 branch_block_stmt_2586/assign_stmt_2931__entry__
      -- CP-element group 1: 	 branch_block_stmt_2586/assign_stmt_2931__exit__
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2586/assign_stmt_2931/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/assign_stmt_2931/$exit
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2702/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_sources/type_cast_2708/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_sources/type_cast_2708/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_sources/type_cast_2708/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_sources/type_cast_2708/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_sources/type_cast_2708/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_sources/type_cast_2708/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2709/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_sources/type_cast_2715/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_sources/type_cast_2715/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_sources/type_cast_2715/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_sources/type_cast_2715/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_sources/type_cast_2715/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_sources/type_cast_2715/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2716/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_sources/type_cast_2722/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_sources/type_cast_2722/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_sources/type_cast_2722/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_sources/type_cast_2722/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_sources/type_cast_2722/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_sources/type_cast_2722/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2723/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2728/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2728/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2728/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2728/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2728/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2728/SplitProtocol/Update/cr
      -- 
    rr_7494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(1), ack => type_cast_2708_inst_req_0); -- 
    cr_7499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(1), ack => type_cast_2708_inst_req_1); -- 
    rr_7517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(1), ack => type_cast_2715_inst_req_0); -- 
    cr_7522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(1), ack => type_cast_2715_inst_req_1); -- 
    rr_7540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(1), ack => type_cast_2722_inst_req_0); -- 
    cr_7545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(1), ack => type_cast_2722_inst_req_1); -- 
    rr_7563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(1), ack => type_cast_2728_inst_req_0); -- 
    cr_7568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(1), ack => type_cast_2728_inst_req_1); -- 
    convTransposeD_CP_6773_elements(1) <= convTransposeD_CP_6773_elements(123);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2588_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2588_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2588_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2588_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2588_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2588_Update/cr
      -- 
    ra_6822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2588_inst_ack_0, ack => convTransposeD_CP_6773_elements(2)); -- 
    cr_6826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(2), ack => RPIPE_Block3_start_2588_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2588_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2588_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2588_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2591_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2591_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2591_Sample/rr
      -- 
    ca_6827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2588_inst_ack_1, ack => convTransposeD_CP_6773_elements(3)); -- 
    rr_6835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(3), ack => RPIPE_Block3_start_2591_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2591_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2591_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2591_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2591_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2591_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2591_Update/cr
      -- 
    ra_6836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2591_inst_ack_0, ack => convTransposeD_CP_6773_elements(4)); -- 
    cr_6840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(4), ack => RPIPE_Block3_start_2591_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2591_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2591_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2591_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2594_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2594_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2594_Sample/rr
      -- 
    ca_6841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2591_inst_ack_1, ack => convTransposeD_CP_6773_elements(5)); -- 
    rr_6849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(5), ack => RPIPE_Block3_start_2594_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2594_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2594_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2594_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2594_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2594_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2594_Update/cr
      -- 
    ra_6850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2594_inst_ack_0, ack => convTransposeD_CP_6773_elements(6)); -- 
    cr_6854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(6), ack => RPIPE_Block3_start_2594_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2594_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2594_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2594_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2597_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2597_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2597_Sample/rr
      -- 
    ca_6855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2594_inst_ack_1, ack => convTransposeD_CP_6773_elements(7)); -- 
    rr_6863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(7), ack => RPIPE_Block3_start_2597_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2597_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2597_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2597_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2597_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2597_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2597_Update/cr
      -- 
    ra_6864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2597_inst_ack_0, ack => convTransposeD_CP_6773_elements(8)); -- 
    cr_6868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(8), ack => RPIPE_Block3_start_2597_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2597_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2597_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2597_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2600_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2600_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2600_Sample/rr
      -- 
    ca_6869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2597_inst_ack_1, ack => convTransposeD_CP_6773_elements(9)); -- 
    rr_6877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(9), ack => RPIPE_Block3_start_2600_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2600_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2600_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2600_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2600_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2600_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2600_Update/cr
      -- 
    ra_6878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2600_inst_ack_0, ack => convTransposeD_CP_6773_elements(10)); -- 
    cr_6882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(10), ack => RPIPE_Block3_start_2600_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2600_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2600_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2600_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2603_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2603_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2603_Sample/rr
      -- 
    ca_6883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2600_inst_ack_1, ack => convTransposeD_CP_6773_elements(11)); -- 
    rr_6891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(11), ack => RPIPE_Block3_start_2603_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2603_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2603_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2603_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2603_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2603_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2603_Update/cr
      -- 
    ra_6892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2603_inst_ack_0, ack => convTransposeD_CP_6773_elements(12)); -- 
    cr_6896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(12), ack => RPIPE_Block3_start_2603_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2603_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2603_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2603_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2606_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2606_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2606_Sample/rr
      -- 
    ca_6897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2603_inst_ack_1, ack => convTransposeD_CP_6773_elements(13)); -- 
    rr_6905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(13), ack => RPIPE_Block3_start_2606_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2606_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2606_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2606_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2606_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2606_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2606_Update/cr
      -- 
    ra_6906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2606_inst_ack_0, ack => convTransposeD_CP_6773_elements(14)); -- 
    cr_6910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(14), ack => RPIPE_Block3_start_2606_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2606_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2606_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2606_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2609_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2609_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2609_Sample/rr
      -- 
    ca_6911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2606_inst_ack_1, ack => convTransposeD_CP_6773_elements(15)); -- 
    rr_6919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(15), ack => RPIPE_Block3_start_2609_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2609_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2609_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2609_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2609_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2609_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2609_Update/cr
      -- 
    ra_6920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2609_inst_ack_0, ack => convTransposeD_CP_6773_elements(16)); -- 
    cr_6924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(16), ack => RPIPE_Block3_start_2609_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2609_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2609_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2609_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2612_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2612_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2612_Sample/rr
      -- 
    ca_6925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2609_inst_ack_1, ack => convTransposeD_CP_6773_elements(17)); -- 
    rr_6933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(17), ack => RPIPE_Block3_start_2612_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2612_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2612_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2612_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2612_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2612_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2612_Update/cr
      -- 
    ra_6934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2612_inst_ack_0, ack => convTransposeD_CP_6773_elements(18)); -- 
    cr_6938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(18), ack => RPIPE_Block3_start_2612_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2612_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2612_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2612_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2615_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2615_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2615_Sample/rr
      -- 
    ca_6939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2612_inst_ack_1, ack => convTransposeD_CP_6773_elements(19)); -- 
    rr_6947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(19), ack => RPIPE_Block3_start_2615_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2615_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2615_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2615_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2615_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2615_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2615_Update/cr
      -- 
    ra_6948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2615_inst_ack_0, ack => convTransposeD_CP_6773_elements(20)); -- 
    cr_6952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(20), ack => RPIPE_Block3_start_2615_inst_req_1); -- 
    -- CP-element group 21:  fork  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (9) 
      -- CP-element group 21: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2628_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2628_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2628_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2615_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2615_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2615_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2619_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2619_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2619_Sample/rr
      -- 
    ca_6953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2615_inst_ack_1, ack => convTransposeD_CP_6773_elements(21)); -- 
    rr_6961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(21), ack => type_cast_2619_inst_req_0); -- 
    rr_6975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(21), ack => RPIPE_Block3_start_2628_inst_req_0); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2619_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2619_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2619_Sample/ra
      -- 
    ra_6962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2619_inst_ack_0, ack => convTransposeD_CP_6773_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	0 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2619_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2619_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2619_update_completed_
      -- 
    ca_6967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2619_inst_ack_1, ack => convTransposeD_CP_6773_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2628_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2628_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2628_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2628_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2628_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2628_update_start_
      -- 
    ra_6976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2628_inst_ack_0, ack => convTransposeD_CP_6773_elements(24)); -- 
    cr_6980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(24), ack => RPIPE_Block3_start_2628_inst_req_1); -- 
    -- CP-element group 25:  fork  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: 	28 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2632_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2640_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2640_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2632_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2640_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2628_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2628_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2632_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2628_update_completed_
      -- 
    ca_6981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2628_inst_ack_1, ack => convTransposeD_CP_6773_elements(25)); -- 
    rr_6989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(25), ack => type_cast_2632_inst_req_0); -- 
    rr_7003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(25), ack => RPIPE_Block3_start_2640_inst_req_0); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2632_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2632_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2632_sample_completed_
      -- 
    ra_6990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2632_inst_ack_0, ack => convTransposeD_CP_6773_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2632_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2632_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/type_cast_2632_update_completed_
      -- 
    ca_6995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2632_inst_ack_1, ack => convTransposeD_CP_6773_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	25 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2640_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2640_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2640_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2640_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2640_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2640_Update/cr
      -- 
    ra_7004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2640_inst_ack_0, ack => convTransposeD_CP_6773_elements(28)); -- 
    cr_7008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(28), ack => RPIPE_Block3_start_2640_inst_req_1); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2643_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2640_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2643_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2640_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2640_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2643_Sample/$entry
      -- 
    ca_7009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2640_inst_ack_1, ack => convTransposeD_CP_6773_elements(29)); -- 
    rr_7017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(29), ack => RPIPE_Block3_start_2643_inst_req_0); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2643_update_start_
      -- CP-element group 30: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2643_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2643_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2643_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2643_Update/cr
      -- CP-element group 30: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2643_Sample/$exit
      -- 
    ra_7018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2643_inst_ack_0, ack => convTransposeD_CP_6773_elements(30)); -- 
    cr_7022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(30), ack => RPIPE_Block3_start_2643_inst_req_1); -- 
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2646_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2643_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2643_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2646_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2646_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2643_update_completed_
      -- 
    ca_7023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2643_inst_ack_1, ack => convTransposeD_CP_6773_elements(31)); -- 
    rr_7031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(31), ack => RPIPE_Block3_start_2646_inst_req_0); -- 
    -- CP-element group 32:  transition  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (6) 
      -- CP-element group 32: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2646_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2646_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2646_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2646_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2646_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2646_Update/$entry
      -- 
    ra_7032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2646_inst_ack_0, ack => convTransposeD_CP_6773_elements(32)); -- 
    cr_7036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(32), ack => RPIPE_Block3_start_2646_inst_req_1); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2646_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2646_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/RPIPE_Block3_start_2646_update_completed_
      -- 
    ca_7037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2646_inst_ack_1, ack => convTransposeD_CP_6773_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  place  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	38 
    -- CP-element group 34: 	39 
    -- CP-element group 34: 	40 
    -- CP-element group 34:  members (22) 
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2694_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2698_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2694_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2694_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2694_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2698_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2690_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2694_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2698_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2690_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2694_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2690_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2698_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2690_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2698_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2698_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2690_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2690_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/$entry
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647__exit__
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699__entry__
      -- CP-element group 34: 	 branch_block_stmt_2586/assign_stmt_2589_to_assign_stmt_2647/$exit
      -- 
    cr_7081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(34), ack => type_cast_2698_inst_req_1); -- 
    rr_7048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(34), ack => type_cast_2690_inst_req_0); -- 
    cr_7067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(34), ack => type_cast_2694_inst_req_1); -- 
    rr_7076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(34), ack => type_cast_2698_inst_req_0); -- 
    rr_7062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(34), ack => type_cast_2694_inst_req_0); -- 
    cr_7053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(34), ack => type_cast_2690_inst_req_1); -- 
    convTransposeD_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(23) & convTransposeD_CP_6773_elements(27) & convTransposeD_CP_6773_elements(33);
      gj_convTransposeD_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2690_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2690_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2690_sample_completed_
      -- 
    ra_7049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2690_inst_ack_0, ack => convTransposeD_CP_6773_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	41 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2690_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2690_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2690_Update/$exit
      -- 
    ca_7054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2690_inst_ack_1, ack => convTransposeD_CP_6773_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2694_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2694_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2694_Sample/ra
      -- 
    ra_7063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2694_inst_ack_0, ack => convTransposeD_CP_6773_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	34 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2694_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2694_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2694_update_completed_
      -- 
    ca_7068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2694_inst_ack_1, ack => convTransposeD_CP_6773_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	34 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2698_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2698_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2698_Sample/$exit
      -- 
    ra_7077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2698_inst_ack_0, ack => convTransposeD_CP_6773_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	34 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2698_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2698_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/type_cast_2698_update_completed_
      -- 
    ca_7082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2698_inst_ack_1, ack => convTransposeD_CP_6773_elements(40)); -- 
    -- CP-element group 41:  join  fork  transition  place  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	36 
    -- CP-element group 41: 	38 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	75 
    -- CP-element group 41: 	76 
    -- CP-element group 41: 	77 
    -- CP-element group 41: 	78 
    -- CP-element group 41: 	79 
    -- CP-element group 41:  members (18) 
      -- CP-element group 41: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699/$exit
      -- CP-element group 41: 	 branch_block_stmt_2586/assign_stmt_2654_to_assign_stmt_2699__exit__
      -- CP-element group 41: 	 branch_block_stmt_2586/entry_whilex_xbody
      -- CP-element group 41: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 41: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2702/$entry
      -- CP-element group 41: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2709/$entry
      -- CP-element group 41: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2716/$entry
      -- CP-element group 41: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2723/$entry
      -- CP-element group 41: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/$entry
      -- CP-element group 41: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/$entry
      -- CP-element group 41: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/$entry
      -- CP-element group 41: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/Sample/rr
      -- CP-element group 41: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/Update/cr
      -- 
    rr_7468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(41), ack => type_cast_2726_inst_req_0); -- 
    cr_7473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(41), ack => type_cast_2726_inst_req_1); -- 
    convTransposeD_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(36) & convTransposeD_CP_6773_elements(38) & convTransposeD_CP_6773_elements(40);
      gj_convTransposeD_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	100 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2763_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2763_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2763_sample_completed_
      -- 
    ra_7094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2763_inst_ack_0, ack => convTransposeD_CP_6773_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	100 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	56 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2763_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2763_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2763_Update/ca
      -- 
    ca_7099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2763_inst_ack_1, ack => convTransposeD_CP_6773_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	100 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2767_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2767_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2767_Sample/ra
      -- 
    ra_7108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2767_inst_ack_0, ack => convTransposeD_CP_6773_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	100 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	56 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2767_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2767_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2767_update_completed_
      -- 
    ca_7113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2767_inst_ack_1, ack => convTransposeD_CP_6773_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	100 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2771_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2771_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2771_Sample/ra
      -- 
    ra_7122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2771_inst_ack_0, ack => convTransposeD_CP_6773_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	100 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	56 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2771_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2771_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2771_update_completed_
      -- 
    ca_7127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2771_inst_ack_1, ack => convTransposeD_CP_6773_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	100 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2801_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2801_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2801_sample_completed_
      -- 
    ra_7136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2801_inst_ack_0, ack => convTransposeD_CP_6773_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	100 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (16) 
      -- CP-element group 49: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2801_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2801_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_final_index_sum_regn_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_index_resized_1
      -- CP-element group 49: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_index_scaled_1
      -- CP-element group 49: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_index_scale_1/scale_rename_req
      -- CP-element group 49: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_index_computed_1
      -- CP-element group 49: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_index_resize_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_index_scale_1/scale_rename_ack
      -- CP-element group 49: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_final_index_sum_regn_Sample/req
      -- CP-element group 49: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_index_resize_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_index_resize_1/index_resize_req
      -- CP-element group 49: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_index_resize_1/index_resize_ack
      -- CP-element group 49: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_index_scale_1/$entry
      -- CP-element group 49: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_index_scale_1/$exit
      -- CP-element group 49: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2801_Update/$exit
      -- 
    ca_7141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2801_inst_ack_1, ack => convTransposeD_CP_6773_elements(49)); -- 
    req_7166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(49), ack => array_obj_ref_2807_index_offset_req_0); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	66 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_final_index_sum_regn_sample_complete
      -- CP-element group 50: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_final_index_sum_regn_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_final_index_sum_regn_Sample/ack
      -- 
    ack_7167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2807_index_offset_ack_0, ack => convTransposeD_CP_6773_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	100 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (11) 
      -- CP-element group 51: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_root_address_calculated
      -- CP-element group 51: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2808_request/$entry
      -- CP-element group 51: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_base_plus_offset/sum_rename_ack
      -- CP-element group 51: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2808_request/req
      -- CP-element group 51: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2808_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_offset_calculated
      -- CP-element group 51: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_final_index_sum_regn_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_final_index_sum_regn_Update/ack
      -- CP-element group 51: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_base_plus_offset/$entry
      -- CP-element group 51: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_base_plus_offset/$exit
      -- CP-element group 51: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_base_plus_offset/sum_rename_req
      -- 
    ack_7172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2807_index_offset_ack_1, ack => convTransposeD_CP_6773_elements(51)); -- 
    req_7181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(51), ack => addr_of_2808_final_reg_req_0); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2808_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2808_request/$exit
      -- CP-element group 52: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2808_request/ack
      -- 
    ack_7182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2808_final_reg_ack_0, ack => convTransposeD_CP_6773_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	100 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (24) 
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2808_complete/ack
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2808_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_base_addr_resize/base_resize_ack
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_base_addr_resize/$entry
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_base_addr_resize/$exit
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2808_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_base_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_base_addr_resize/base_resize_req
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_base_plus_offset/$entry
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_base_plus_offset/$exit
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_word_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_root_address_calculated
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_base_address_resized
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_base_plus_offset/sum_rename_req
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_base_plus_offset/sum_rename_ack
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_word_addrgen/$entry
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_word_addrgen/$exit
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_word_addrgen/root_register_req
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_word_addrgen/root_register_ack
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Sample/word_access_start/word_0/rr
      -- 
    ack_7187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2808_final_reg_ack_1, ack => convTransposeD_CP_6773_elements(53)); -- 
    rr_7220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(53), ack => ptr_deref_2812_load_0_req_0); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Sample/word_access_start/word_0/ra
      -- 
    ra_7221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2812_load_0_ack_0, ack => convTransposeD_CP_6773_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	100 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	61 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Update/word_access_complete/word_0/ca
      -- CP-element group 55: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Update/ptr_deref_2812_Merge/$entry
      -- CP-element group 55: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Update/ptr_deref_2812_Merge/$exit
      -- CP-element group 55: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Update/ptr_deref_2812_Merge/merge_req
      -- CP-element group 55: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Update/ptr_deref_2812_Merge/merge_ack
      -- 
    ca_7232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2812_load_0_ack_1, ack => convTransposeD_CP_6773_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	43 
    -- CP-element group 56: 	45 
    -- CP-element group 56: 	47 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (13) 
      -- CP-element group 56: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_index_scale_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_index_resized_1
      -- CP-element group 56: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_index_scaled_1
      -- CP-element group 56: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_index_computed_1
      -- CP-element group 56: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_index_resize_1/$entry
      -- CP-element group 56: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_index_resize_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_index_resize_1/index_resize_req
      -- CP-element group 56: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_index_resize_1/index_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_index_scale_1/$exit
      -- CP-element group 56: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_index_scale_1/scale_rename_req
      -- CP-element group 56: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_index_scale_1/scale_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_final_index_sum_regn_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_final_index_sum_regn_Sample/req
      -- 
    req_7262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(56), ack => array_obj_ref_2830_index_offset_req_0); -- 
    convTransposeD_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(43) & convTransposeD_CP_6773_elements(45) & convTransposeD_CP_6773_elements(47);
      gj_convTransposeD_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	66 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_final_index_sum_regn_sample_complete
      -- CP-element group 57: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_final_index_sum_regn_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_final_index_sum_regn_Sample/ack
      -- 
    ack_7263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2830_index_offset_ack_0, ack => convTransposeD_CP_6773_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	100 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (11) 
      -- CP-element group 58: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2831_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_root_address_calculated
      -- CP-element group 58: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_offset_calculated
      -- CP-element group 58: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_final_index_sum_regn_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_final_index_sum_regn_Update/ack
      -- CP-element group 58: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_base_plus_offset/$entry
      -- CP-element group 58: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_base_plus_offset/$exit
      -- CP-element group 58: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_base_plus_offset/sum_rename_req
      -- CP-element group 58: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_base_plus_offset/sum_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2831_request/$entry
      -- CP-element group 58: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2831_request/req
      -- 
    ack_7268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2830_index_offset_ack_1, ack => convTransposeD_CP_6773_elements(58)); -- 
    req_7277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(58), ack => addr_of_2831_final_reg_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2831_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2831_request/$exit
      -- CP-element group 59: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2831_request/ack
      -- 
    ack_7278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2831_final_reg_ack_0, ack => convTransposeD_CP_6773_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	100 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (19) 
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2831_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2831_complete/$exit
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2831_complete/ack
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_base_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_word_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_base_address_resized
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_base_addr_resize/$entry
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_base_addr_resize/$exit
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_base_addr_resize/base_resize_req
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_base_addr_resize/base_resize_ack
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_base_plus_offset/sum_rename_ack
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_word_addrgen/$entry
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_word_addrgen/$exit
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_word_addrgen/root_register_req
      -- CP-element group 60: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_word_addrgen/root_register_ack
      -- 
    ack_7283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2831_final_reg_ack_1, ack => convTransposeD_CP_6773_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	55 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (9) 
      -- CP-element group 61: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Sample/ptr_deref_2834_Split/$entry
      -- CP-element group 61: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Sample/ptr_deref_2834_Split/$exit
      -- CP-element group 61: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Sample/ptr_deref_2834_Split/split_req
      -- CP-element group 61: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Sample/ptr_deref_2834_Split/split_ack
      -- CP-element group 61: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Sample/word_access_start/$entry
      -- CP-element group 61: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Sample/word_access_start/word_0/$entry
      -- CP-element group 61: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Sample/word_access_start/word_0/rr
      -- 
    rr_7321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(61), ack => ptr_deref_2834_store_0_req_0); -- 
    convTransposeD_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(55) & convTransposeD_CP_6773_elements(60);
      gj_convTransposeD_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (5) 
      -- CP-element group 62: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Sample/word_access_start/$exit
      -- CP-element group 62: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Sample/word_access_start/word_0/$exit
      -- CP-element group 62: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Sample/word_access_start/word_0/ra
      -- 
    ra_7322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_store_0_ack_0, ack => convTransposeD_CP_6773_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	100 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (5) 
      -- CP-element group 63: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Update/word_access_complete/$exit
      -- CP-element group 63: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Update/word_access_complete/word_0/$exit
      -- CP-element group 63: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Update/word_access_complete/word_0/ca
      -- 
    ca_7333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_store_0_ack_1, ack => convTransposeD_CP_6773_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	100 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2839_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2839_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2839_Sample/ra
      -- 
    ra_7342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2839_inst_ack_0, ack => convTransposeD_CP_6773_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	100 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2839_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2839_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2839_Update/ca
      -- 
    ca_7347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2839_inst_ack_1, ack => convTransposeD_CP_6773_elements(65)); -- 
    -- CP-element group 66:  branch  join  transition  place  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	50 
    -- CP-element group 66: 	57 
    -- CP-element group 66: 	63 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (10) 
      -- CP-element group 66: 	 branch_block_stmt_2586/R_cmp_2853_place
      -- CP-element group 66: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/$exit
      -- CP-element group 66: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851__exit__
      -- CP-element group 66: 	 branch_block_stmt_2586/if_stmt_2852__entry__
      -- CP-element group 66: 	 branch_block_stmt_2586/if_stmt_2852_dead_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2586/if_stmt_2852_eval_test/$entry
      -- CP-element group 66: 	 branch_block_stmt_2586/if_stmt_2852_eval_test/$exit
      -- CP-element group 66: 	 branch_block_stmt_2586/if_stmt_2852_eval_test/branch_req
      -- CP-element group 66: 	 branch_block_stmt_2586/if_stmt_2852_if_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2586/if_stmt_2852_else_link/$entry
      -- 
    branch_req_7355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(66), ack => if_stmt_2852_branch_req_0); -- 
    convTransposeD_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(50) & convTransposeD_CP_6773_elements(57) & convTransposeD_CP_6773_elements(63) & convTransposeD_CP_6773_elements(65);
      gj_convTransposeD_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	109 
    -- CP-element group 67: 	110 
    -- CP-element group 67: 	112 
    -- CP-element group 67: 	113 
    -- CP-element group 67: 	115 
    -- CP-element group 67: 	116 
    -- CP-element group 67:  members (40) 
      -- CP-element group 67: 	 branch_block_stmt_2586/whilex_xbody_ifx_xthen
      -- CP-element group 67: 	 branch_block_stmt_2586/merge_stmt_2858__exit__
      -- CP-element group 67: 	 branch_block_stmt_2586/assign_stmt_2864__entry__
      -- CP-element group 67: 	 branch_block_stmt_2586/assign_stmt_2864__exit__
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132
      -- CP-element group 67: 	 branch_block_stmt_2586/if_stmt_2852_if_link/$exit
      -- CP-element group 67: 	 branch_block_stmt_2586/if_stmt_2852_if_link/if_choice_transition
      -- CP-element group 67: 	 branch_block_stmt_2586/assign_stmt_2864/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/assign_stmt_2864/$exit
      -- CP-element group 67: 	 branch_block_stmt_2586/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_2586/merge_stmt_2858_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_2586/merge_stmt_2858_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/merge_stmt_2858_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_2586/merge_stmt_2858_PhiAck/dummy
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2906/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_sources/type_cast_2909/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_sources/type_cast_2909/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_sources/type_cast_2909/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_sources/type_cast_2909/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_sources/type_cast_2909/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_sources/type_cast_2909/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/Update/cr
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2919/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2922/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2922/SplitProtocol/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2922/SplitProtocol/Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2922/SplitProtocol/Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2922/SplitProtocol/Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2922/SplitProtocol/Update/cr
      -- 
    if_choice_transition_7360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2852_branch_ack_1, ack => convTransposeD_CP_6773_elements(67)); -- 
    rr_7678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(67), ack => type_cast_2909_inst_req_0); -- 
    cr_7683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(67), ack => type_cast_2909_inst_req_1); -- 
    rr_7701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(67), ack => type_cast_2916_inst_req_0); -- 
    cr_7706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(67), ack => type_cast_2916_inst_req_1); -- 
    rr_7724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(67), ack => type_cast_2922_inst_req_0); -- 
    cr_7729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(67), ack => type_cast_2922_inst_req_1); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (18) 
      -- CP-element group 68: 	 branch_block_stmt_2586/whilex_xbody_ifx_xelse
      -- CP-element group 68: 	 branch_block_stmt_2586/merge_stmt_2866__exit__
      -- CP-element group 68: 	 branch_block_stmt_2586/assign_stmt_2872_to_assign_stmt_2898__entry__
      -- CP-element group 68: 	 branch_block_stmt_2586/if_stmt_2852_else_link/$exit
      -- CP-element group 68: 	 branch_block_stmt_2586/if_stmt_2852_else_link/else_choice_transition
      -- CP-element group 68: 	 branch_block_stmt_2586/assign_stmt_2872_to_assign_stmt_2898/$entry
      -- CP-element group 68: 	 branch_block_stmt_2586/assign_stmt_2872_to_assign_stmt_2898/type_cast_2880_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_2586/assign_stmt_2872_to_assign_stmt_2898/type_cast_2880_update_start_
      -- CP-element group 68: 	 branch_block_stmt_2586/assign_stmt_2872_to_assign_stmt_2898/type_cast_2880_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2586/assign_stmt_2872_to_assign_stmt_2898/type_cast_2880_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2586/assign_stmt_2872_to_assign_stmt_2898/type_cast_2880_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2586/assign_stmt_2872_to_assign_stmt_2898/type_cast_2880_Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2586/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2586/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_2586/merge_stmt_2866_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_2586/merge_stmt_2866_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_2586/merge_stmt_2866_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_2586/merge_stmt_2866_PhiAck/dummy
      -- 
    else_choice_transition_7364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2852_branch_ack_0, ack => convTransposeD_CP_6773_elements(68)); -- 
    rr_7380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(68), ack => type_cast_2880_inst_req_0); -- 
    cr_7385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(68), ack => type_cast_2880_inst_req_1); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2586/assign_stmt_2872_to_assign_stmt_2898/type_cast_2880_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2586/assign_stmt_2872_to_assign_stmt_2898/type_cast_2880_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2586/assign_stmt_2872_to_assign_stmt_2898/type_cast_2880_Sample/ra
      -- 
    ra_7381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2880_inst_ack_0, ack => convTransposeD_CP_6773_elements(69)); -- 
    -- CP-element group 70:  branch  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (13) 
      -- CP-element group 70: 	 branch_block_stmt_2586/assign_stmt_2872_to_assign_stmt_2898__exit__
      -- CP-element group 70: 	 branch_block_stmt_2586/if_stmt_2899__entry__
      -- CP-element group 70: 	 branch_block_stmt_2586/assign_stmt_2872_to_assign_stmt_2898/$exit
      -- CP-element group 70: 	 branch_block_stmt_2586/assign_stmt_2872_to_assign_stmt_2898/type_cast_2880_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2586/assign_stmt_2872_to_assign_stmt_2898/type_cast_2880_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2586/assign_stmt_2872_to_assign_stmt_2898/type_cast_2880_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_2586/if_stmt_2899_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2586/if_stmt_2899_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_2586/if_stmt_2899_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_2586/if_stmt_2899_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_2586/R_cmp121_2900_place
      -- CP-element group 70: 	 branch_block_stmt_2586/if_stmt_2899_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2586/if_stmt_2899_else_link/$entry
      -- 
    ca_7386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2880_inst_ack_1, ack => convTransposeD_CP_6773_elements(70)); -- 
    branch_req_7394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(70), ack => if_stmt_2899_branch_req_0); -- 
    -- CP-element group 71:  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (15) 
      -- CP-element group 71: 	 branch_block_stmt_2586/merge_stmt_2933__exit__
      -- CP-element group 71: 	 branch_block_stmt_2586/assign_stmt_2938__entry__
      -- CP-element group 71: 	 branch_block_stmt_2586/if_stmt_2899_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_2586/if_stmt_2899_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_2586/ifx_xelse_whilex_xend
      -- CP-element group 71: 	 branch_block_stmt_2586/assign_stmt_2938/$entry
      -- CP-element group 71: 	 branch_block_stmt_2586/assign_stmt_2938/WPIPE_Block3_done_2935_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2586/assign_stmt_2938/WPIPE_Block3_done_2935_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2586/assign_stmt_2938/WPIPE_Block3_done_2935_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_2586/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_2586/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_2586/merge_stmt_2933_PhiReqMerge
      -- CP-element group 71: 	 branch_block_stmt_2586/merge_stmt_2933_PhiAck/$entry
      -- CP-element group 71: 	 branch_block_stmt_2586/merge_stmt_2933_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_2586/merge_stmt_2933_PhiAck/dummy
      -- 
    if_choice_transition_7399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2899_branch_ack_1, ack => convTransposeD_CP_6773_elements(71)); -- 
    req_7419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(71), ack => WPIPE_Block3_done_2935_inst_req_0); -- 
    -- CP-element group 72:  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	101 
    -- CP-element group 72: 	102 
    -- CP-element group 72: 	103 
    -- CP-element group 72: 	105 
    -- CP-element group 72: 	106 
    -- CP-element group 72:  members (22) 
      -- CP-element group 72: 	 branch_block_stmt_2586/if_stmt_2899_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_2586/if_stmt_2899_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2906/$entry
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/$entry
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/$entry
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2919/$entry
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2924/$entry
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2924/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2924/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2924/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2924/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2924/SplitProtocol/Update/cr
      -- 
    else_choice_transition_7403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2899_branch_ack_0, ack => convTransposeD_CP_6773_elements(72)); -- 
    rr_7629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(72), ack => type_cast_2918_inst_req_0); -- 
    cr_7634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(72), ack => type_cast_2918_inst_req_1); -- 
    rr_7652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(72), ack => type_cast_2924_inst_req_0); -- 
    cr_7657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(72), ack => type_cast_2924_inst_req_1); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_2586/assign_stmt_2938/WPIPE_Block3_done_2935_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2586/assign_stmt_2938/WPIPE_Block3_done_2935_update_start_
      -- CP-element group 73: 	 branch_block_stmt_2586/assign_stmt_2938/WPIPE_Block3_done_2935_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2586/assign_stmt_2938/WPIPE_Block3_done_2935_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_2586/assign_stmt_2938/WPIPE_Block3_done_2935_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_2586/assign_stmt_2938/WPIPE_Block3_done_2935_Update/req
      -- 
    ack_7420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2935_inst_ack_0, ack => convTransposeD_CP_6773_elements(73)); -- 
    req_7424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(73), ack => WPIPE_Block3_done_2935_inst_req_1); -- 
    -- CP-element group 74:  transition  place  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (16) 
      -- CP-element group 74: 	 $exit
      -- CP-element group 74: 	 branch_block_stmt_2586/$exit
      -- CP-element group 74: 	 branch_block_stmt_2586/branch_block_stmt_2586__exit__
      -- CP-element group 74: 	 branch_block_stmt_2586/assign_stmt_2938__exit__
      -- CP-element group 74: 	 branch_block_stmt_2586/return__
      -- CP-element group 74: 	 branch_block_stmt_2586/merge_stmt_2940__exit__
      -- CP-element group 74: 	 branch_block_stmt_2586/assign_stmt_2938/$exit
      -- CP-element group 74: 	 branch_block_stmt_2586/assign_stmt_2938/WPIPE_Block3_done_2935_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2586/assign_stmt_2938/WPIPE_Block3_done_2935_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2586/assign_stmt_2938/WPIPE_Block3_done_2935_Update/ack
      -- CP-element group 74: 	 branch_block_stmt_2586/return___PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_2586/return___PhiReq/$exit
      -- CP-element group 74: 	 branch_block_stmt_2586/merge_stmt_2940_PhiReqMerge
      -- CP-element group 74: 	 branch_block_stmt_2586/merge_stmt_2940_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_2586/merge_stmt_2940_PhiAck/$exit
      -- CP-element group 74: 	 branch_block_stmt_2586/merge_stmt_2940_PhiAck/dummy
      -- 
    ack_7425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2935_inst_ack_1, ack => convTransposeD_CP_6773_elements(74)); -- 
    -- CP-element group 75:  transition  output  delay-element  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	41 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	81 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2702/$exit
      -- CP-element group 75: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_sources/type_cast_2706_konst_delay_trans
      -- CP-element group 75: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_req
      -- 
    phi_stmt_2702_req_7436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2702_req_7436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(75), ack => phi_stmt_2702_req_0); -- 
    -- Element group convTransposeD_CP_6773_elements(75) is a control-delay.
    cp_element_75_delay: control_delay_element  generic map(name => " 75_delay", delay_value => 1)  port map(req => convTransposeD_CP_6773_elements(41), ack => convTransposeD_CP_6773_elements(75), clk => clk, reset =>reset);
    -- CP-element group 76:  transition  output  delay-element  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	41 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	81 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2709/$exit
      -- CP-element group 76: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_sources/type_cast_2713_konst_delay_trans
      -- CP-element group 76: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_req
      -- 
    phi_stmt_2709_req_7444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2709_req_7444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(76), ack => phi_stmt_2709_req_0); -- 
    -- Element group convTransposeD_CP_6773_elements(76) is a control-delay.
    cp_element_76_delay: control_delay_element  generic map(name => " 76_delay", delay_value => 1)  port map(req => convTransposeD_CP_6773_elements(41), ack => convTransposeD_CP_6773_elements(76), clk => clk, reset =>reset);
    -- CP-element group 77:  transition  output  delay-element  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	41 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2716/$exit
      -- CP-element group 77: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_sources/type_cast_2720_konst_delay_trans
      -- CP-element group 77: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_req
      -- 
    phi_stmt_2716_req_7452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2716_req_7452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(77), ack => phi_stmt_2716_req_0); -- 
    -- Element group convTransposeD_CP_6773_elements(77) is a control-delay.
    cp_element_77_delay: control_delay_element  generic map(name => " 77_delay", delay_value => 1)  port map(req => convTransposeD_CP_6773_elements(41), ack => convTransposeD_CP_6773_elements(77), clk => clk, reset =>reset);
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	41 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/Sample/ra
      -- 
    ra_7469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2726_inst_ack_0, ack => convTransposeD_CP_6773_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	41 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/Update/ca
      -- 
    ca_7474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2726_inst_ack_1, ack => convTransposeD_CP_6773_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2723/$exit
      -- CP-element group 80: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/$exit
      -- CP-element group 80: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2726/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_req
      -- 
    phi_stmt_2723_req_7475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2723_req_7475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(80), ack => phi_stmt_2723_req_0); -- 
    convTransposeD_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(78) & convTransposeD_CP_6773_elements(79);
      gj_convTransposeD_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: 	76 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	95 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2586/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(75) & convTransposeD_CP_6773_elements(76) & convTransposeD_CP_6773_elements(77) & convTransposeD_CP_6773_elements(80);
      gj_convTransposeD_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	1 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_sources/type_cast_2708/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_sources/type_cast_2708/SplitProtocol/Sample/ra
      -- 
    ra_7495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2708_inst_ack_0, ack => convTransposeD_CP_6773_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	1 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_sources/type_cast_2708/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_sources/type_cast_2708/SplitProtocol/Update/ca
      -- 
    ca_7500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2708_inst_ack_1, ack => convTransposeD_CP_6773_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	94 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2702/$exit
      -- CP-element group 84: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_sources/type_cast_2708/$exit
      -- CP-element group 84: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_sources/type_cast_2708/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2702/phi_stmt_2702_req
      -- 
    phi_stmt_2702_req_7501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2702_req_7501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(84), ack => phi_stmt_2702_req_1); -- 
    convTransposeD_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(82) & convTransposeD_CP_6773_elements(83);
      gj_convTransposeD_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	1 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_sources/type_cast_2715/SplitProtocol/Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_sources/type_cast_2715/SplitProtocol/Sample/ra
      -- 
    ra_7518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2715_inst_ack_0, ack => convTransposeD_CP_6773_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	1 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_sources/type_cast_2715/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_sources/type_cast_2715/SplitProtocol/Update/ca
      -- 
    ca_7523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2715_inst_ack_1, ack => convTransposeD_CP_6773_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	94 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2709/$exit
      -- CP-element group 87: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_sources/type_cast_2715/$exit
      -- CP-element group 87: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_sources/type_cast_2715/SplitProtocol/$exit
      -- CP-element group 87: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2709/phi_stmt_2709_req
      -- 
    phi_stmt_2709_req_7524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2709_req_7524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(87), ack => phi_stmt_2709_req_1); -- 
    convTransposeD_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(85) & convTransposeD_CP_6773_elements(86);
      gj_convTransposeD_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	1 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_sources/type_cast_2722/SplitProtocol/Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_sources/type_cast_2722/SplitProtocol/Sample/ra
      -- 
    ra_7541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2722_inst_ack_0, ack => convTransposeD_CP_6773_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	1 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_sources/type_cast_2722/SplitProtocol/Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_sources/type_cast_2722/SplitProtocol/Update/ca
      -- 
    ca_7546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2722_inst_ack_1, ack => convTransposeD_CP_6773_elements(89)); -- 
    -- CP-element group 90:  join  transition  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	94 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2716/$exit
      -- CP-element group 90: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_sources/$exit
      -- CP-element group 90: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_sources/type_cast_2722/$exit
      -- CP-element group 90: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_sources/type_cast_2722/SplitProtocol/$exit
      -- CP-element group 90: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2716/phi_stmt_2716_req
      -- 
    phi_stmt_2716_req_7547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2716_req_7547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(90), ack => phi_stmt_2716_req_1); -- 
    convTransposeD_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(88) & convTransposeD_CP_6773_elements(89);
      gj_convTransposeD_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	1 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2728/SplitProtocol/Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2728/SplitProtocol/Sample/ra
      -- 
    ra_7564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2728_inst_ack_0, ack => convTransposeD_CP_6773_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	1 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (2) 
      -- CP-element group 92: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2728/SplitProtocol/Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2728/SplitProtocol/Update/ca
      -- 
    ca_7569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2728_inst_ack_1, ack => convTransposeD_CP_6773_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2723/$exit
      -- CP-element group 93: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2728/$exit
      -- CP-element group 93: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_sources/type_cast_2728/SplitProtocol/$exit
      -- CP-element group 93: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/phi_stmt_2723/phi_stmt_2723_req
      -- 
    phi_stmt_2723_req_7570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2723_req_7570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(93), ack => phi_stmt_2723_req_1); -- 
    convTransposeD_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(91) & convTransposeD_CP_6773_elements(92);
      gj_convTransposeD_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	84 
    -- CP-element group 94: 	87 
    -- CP-element group 94: 	90 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_2586/ifx_xend132_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(84) & convTransposeD_CP_6773_elements(87) & convTransposeD_CP_6773_elements(90) & convTransposeD_CP_6773_elements(93);
      gj_convTransposeD_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  merge  fork  transition  place  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	81 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	97 
    -- CP-element group 95: 	98 
    -- CP-element group 95: 	99 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2586/merge_stmt_2701_PhiReqMerge
      -- CP-element group 95: 	 branch_block_stmt_2586/merge_stmt_2701_PhiAck/$entry
      -- 
    convTransposeD_CP_6773_elements(95) <= OrReduce(convTransposeD_CP_6773_elements(81) & convTransposeD_CP_6773_elements(94));
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	100 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_2586/merge_stmt_2701_PhiAck/phi_stmt_2702_ack
      -- 
    phi_stmt_2702_ack_7575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2702_ack_0, ack => convTransposeD_CP_6773_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	100 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_2586/merge_stmt_2701_PhiAck/phi_stmt_2709_ack
      -- 
    phi_stmt_2709_ack_7576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2709_ack_0, ack => convTransposeD_CP_6773_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2586/merge_stmt_2701_PhiAck/phi_stmt_2716_ack
      -- 
    phi_stmt_2716_ack_7577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2716_ack_0, ack => convTransposeD_CP_6773_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	95 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_2586/merge_stmt_2701_PhiAck/phi_stmt_2723_ack
      -- 
    phi_stmt_2723_ack_7578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2723_ack_0, ack => convTransposeD_CP_6773_elements(99)); -- 
    -- CP-element group 100:  join  fork  transition  place  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	96 
    -- CP-element group 100: 	97 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	42 
    -- CP-element group 100: 	43 
    -- CP-element group 100: 	44 
    -- CP-element group 100: 	45 
    -- CP-element group 100: 	46 
    -- CP-element group 100: 	47 
    -- CP-element group 100: 	48 
    -- CP-element group 100: 	49 
    -- CP-element group 100: 	51 
    -- CP-element group 100: 	53 
    -- CP-element group 100: 	55 
    -- CP-element group 100: 	58 
    -- CP-element group 100: 	60 
    -- CP-element group 100: 	63 
    -- CP-element group 100: 	64 
    -- CP-element group 100: 	65 
    -- CP-element group 100:  members (56) 
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2763_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2801_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2767_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2801_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2808_complete/req
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2808_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2763_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2801_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2763_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2808_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2767_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2771_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2763_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_final_index_sum_regn_update_start
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2767_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2771_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2767_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2801_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2771_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2801_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2771_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_final_index_sum_regn_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2763_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2771_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2807_final_index_sum_regn_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2767_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2767_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2801_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2771_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2763_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2586/merge_stmt_2701__exit__
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851__entry__
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Update/word_access_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Update/word_access_complete/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2812_Update/word_access_complete/word_0/cr
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2831_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_final_index_sum_regn_update_start
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_final_index_sum_regn_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/array_obj_ref_2830_final_index_sum_regn_Update/req
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2831_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/addr_of_2831_complete/req
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Update/word_access_complete/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Update/word_access_complete/word_0/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/ptr_deref_2834_Update/word_access_complete/word_0/cr
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2839_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2839_update_start_
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2839_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2839_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2839_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_2586/assign_stmt_2735_to_assign_stmt_2851/type_cast_2839_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_2586/merge_stmt_2701_PhiAck/$exit
      -- 
    cr_7140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2801_inst_req_1); -- 
    req_7186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => addr_of_2808_final_reg_req_1); -- 
    rr_7135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2801_inst_req_0); -- 
    rr_7093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2763_inst_req_0); -- 
    cr_7112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2767_inst_req_1); -- 
    rr_7107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2767_inst_req_0); -- 
    rr_7121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2771_inst_req_0); -- 
    cr_7126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2771_inst_req_1); -- 
    req_7171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => array_obj_ref_2807_index_offset_req_1); -- 
    cr_7098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2763_inst_req_1); -- 
    cr_7231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => ptr_deref_2812_load_0_req_1); -- 
    req_7267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => array_obj_ref_2830_index_offset_req_1); -- 
    req_7282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => addr_of_2831_final_reg_req_1); -- 
    cr_7332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => ptr_deref_2834_store_0_req_1); -- 
    rr_7341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2839_inst_req_0); -- 
    cr_7346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(100), ack => type_cast_2839_inst_req_1); -- 
    convTransposeD_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(96) & convTransposeD_CP_6773_elements(97) & convTransposeD_CP_6773_elements(98) & convTransposeD_CP_6773_elements(99);
      gj_convTransposeD_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  output  delay-element  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	72 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	108 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2906/$exit
      -- CP-element group 101: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_sources/type_cast_2912_konst_delay_trans
      -- CP-element group 101: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_req
      -- 
    phi_stmt_2906_req_7613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2906_req_7613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(101), ack => phi_stmt_2906_req_1); -- 
    -- Element group convTransposeD_CP_6773_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => convTransposeD_CP_6773_elements(72), ack => convTransposeD_CP_6773_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	72 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/Sample/ra
      -- 
    ra_7630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2918_inst_ack_0, ack => convTransposeD_CP_6773_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	72 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/Update/ca
      -- 
    ca_7635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2918_inst_ack_1, ack => convTransposeD_CP_6773_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/$exit
      -- CP-element group 104: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/$exit
      -- CP-element group 104: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2918/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_req
      -- 
    phi_stmt_2913_req_7636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2913_req_7636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(104), ack => phi_stmt_2913_req_1); -- 
    convTransposeD_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(102) & convTransposeD_CP_6773_elements(103);
      gj_convTransposeD_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	72 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2924/SplitProtocol/Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2924/SplitProtocol/Sample/ra
      -- 
    ra_7653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2924_inst_ack_0, ack => convTransposeD_CP_6773_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	72 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2924/SplitProtocol/Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2924/SplitProtocol/Update/ca
      -- 
    ca_7658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2924_inst_ack_1, ack => convTransposeD_CP_6773_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2919/$exit
      -- CP-element group 107: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2924/$exit
      -- CP-element group 107: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2924/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_req
      -- 
    phi_stmt_2919_req_7659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2919_req_7659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(107), ack => phi_stmt_2919_req_1); -- 
    convTransposeD_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(105) & convTransposeD_CP_6773_elements(106);
      gj_convTransposeD_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	101 
    -- CP-element group 108: 	104 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	119 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_2586/ifx_xelse_ifx_xend132_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(101) & convTransposeD_CP_6773_elements(104) & convTransposeD_CP_6773_elements(107);
      gj_convTransposeD_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	67 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_sources/type_cast_2909/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_sources/type_cast_2909/SplitProtocol/Sample/ra
      -- 
    ra_7679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2909_inst_ack_0, ack => convTransposeD_CP_6773_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	67 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_sources/type_cast_2909/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_sources/type_cast_2909/SplitProtocol/Update/ca
      -- 
    ca_7684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2909_inst_ack_1, ack => convTransposeD_CP_6773_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	118 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2906/$exit
      -- CP-element group 111: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_sources/type_cast_2909/$exit
      -- CP-element group 111: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_sources/type_cast_2909/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2906/phi_stmt_2906_req
      -- 
    phi_stmt_2906_req_7685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2906_req_7685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(111), ack => phi_stmt_2906_req_0); -- 
    convTransposeD_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(109) & convTransposeD_CP_6773_elements(110);
      gj_convTransposeD_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	67 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/Sample/ra
      -- 
    ra_7702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2916_inst_ack_0, ack => convTransposeD_CP_6773_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	67 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/Update/ca
      -- 
    ca_7707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2916_inst_ack_1, ack => convTransposeD_CP_6773_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	118 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/$exit
      -- CP-element group 114: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/$exit
      -- CP-element group 114: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/$exit
      -- CP-element group 114: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_sources/type_cast_2916/SplitProtocol/$exit
      -- CP-element group 114: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2913/phi_stmt_2913_req
      -- 
    phi_stmt_2913_req_7708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2913_req_7708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(114), ack => phi_stmt_2913_req_0); -- 
    convTransposeD_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(112) & convTransposeD_CP_6773_elements(113);
      gj_convTransposeD_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	67 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2922/SplitProtocol/Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2922/SplitProtocol/Sample/ra
      -- 
    ra_7725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2922_inst_ack_0, ack => convTransposeD_CP_6773_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	67 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2922/SplitProtocol/Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2922/SplitProtocol/Update/ca
      -- 
    ca_7730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2922_inst_ack_1, ack => convTransposeD_CP_6773_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2919/$exit
      -- CP-element group 117: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/$exit
      -- CP-element group 117: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2922/$exit
      -- CP-element group 117: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_sources/type_cast_2922/SplitProtocol/$exit
      -- CP-element group 117: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/phi_stmt_2919/phi_stmt_2919_req
      -- 
    phi_stmt_2919_req_7731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2919_req_7731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6773_elements(117), ack => phi_stmt_2919_req_0); -- 
    convTransposeD_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(115) & convTransposeD_CP_6773_elements(116);
      gj_convTransposeD_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	111 
    -- CP-element group 118: 	114 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_2586/ifx_xthen_ifx_xend132_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(111) & convTransposeD_CP_6773_elements(114) & convTransposeD_CP_6773_elements(117);
      gj_convTransposeD_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  merge  fork  transition  place  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	108 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119: 	121 
    -- CP-element group 119: 	122 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2586/merge_stmt_2905_PhiReqMerge
      -- CP-element group 119: 	 branch_block_stmt_2586/merge_stmt_2905_PhiAck/$entry
      -- 
    convTransposeD_CP_6773_elements(119) <= OrReduce(convTransposeD_CP_6773_elements(108) & convTransposeD_CP_6773_elements(118));
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	123 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_2586/merge_stmt_2905_PhiAck/phi_stmt_2906_ack
      -- 
    phi_stmt_2906_ack_7736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2906_ack_0, ack => convTransposeD_CP_6773_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_2586/merge_stmt_2905_PhiAck/phi_stmt_2913_ack
      -- 
    phi_stmt_2913_ack_7737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2913_ack_0, ack => convTransposeD_CP_6773_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	119 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_2586/merge_stmt_2905_PhiAck/phi_stmt_2919_ack
      -- 
    phi_stmt_2919_ack_7738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2919_ack_0, ack => convTransposeD_CP_6773_elements(122)); -- 
    -- CP-element group 123:  join  transition  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	120 
    -- CP-element group 123: 	121 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	1 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_2586/merge_stmt_2905_PhiAck/$exit
      -- 
    convTransposeD_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6773_elements(120) & convTransposeD_CP_6773_elements(121) & convTransposeD_CP_6773_elements(122);
      gj_convTransposeD_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6773_elements(123), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom91_2829_resized : std_logic_vector(13 downto 0);
    signal R_idxprom91_2829_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2806_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2806_scaled : std_logic_vector(13 downto 0);
    signal add103_2864 : std_logic_vector(15 downto 0);
    signal add32_2665 : std_logic_vector(15 downto 0);
    signal add50_2671 : std_logic_vector(15 downto 0);
    signal add63_2682 : std_logic_vector(15 downto 0);
    signal add82_2782 : std_logic_vector(63 downto 0);
    signal add84_2792 : std_logic_vector(63 downto 0);
    signal add96_2846 : std_logic_vector(31 downto 0);
    signal add_2638 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2740 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2807_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2807_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2807_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2807_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2807_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2807_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2830_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2830_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2830_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2830_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2830_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2830_root_address : std_logic_vector(13 downto 0);
    signal arrayidx87_2809 : std_logic_vector(31 downto 0);
    signal arrayidx92_2832 : std_logic_vector(31 downto 0);
    signal call11_2607 : std_logic_vector(15 downto 0);
    signal call13_2610 : std_logic_vector(15 downto 0);
    signal call14_2613 : std_logic_vector(15 downto 0);
    signal call15_2616 : std_logic_vector(15 downto 0);
    signal call16_2629 : std_logic_vector(15 downto 0);
    signal call18_2641 : std_logic_vector(15 downto 0);
    signal call1_2592 : std_logic_vector(15 downto 0);
    signal call20_2644 : std_logic_vector(15 downto 0);
    signal call22_2647 : std_logic_vector(15 downto 0);
    signal call3_2595 : std_logic_vector(15 downto 0);
    signal call5_2598 : std_logic_vector(15 downto 0);
    signal call7_2601 : std_logic_vector(15 downto 0);
    signal call9_2604 : std_logic_vector(15 downto 0);
    signal call_2589 : std_logic_vector(15 downto 0);
    signal cmp111_2877 : std_logic_vector(0 downto 0);
    signal cmp121_2898 : std_logic_vector(0 downto 0);
    signal cmp_2851 : std_logic_vector(0 downto 0);
    signal conv17_2633 : std_logic_vector(31 downto 0);
    signal conv70_2764 : std_logic_vector(63 downto 0);
    signal conv73_2691 : std_logic_vector(63 downto 0);
    signal conv75_2768 : std_logic_vector(63 downto 0);
    signal conv78_2695 : std_logic_vector(63 downto 0);
    signal conv80_2772 : std_logic_vector(63 downto 0);
    signal conv95_2840 : std_logic_vector(31 downto 0);
    signal conv99_2699 : std_logic_vector(31 downto 0);
    signal conv_2620 : std_logic_vector(31 downto 0);
    signal idxprom91_2825 : std_logic_vector(63 downto 0);
    signal idxprom_2802 : std_logic_vector(63 downto 0);
    signal inc115_2881 : std_logic_vector(15 downto 0);
    signal inc115x_xinput_dim0x_x2_2886 : std_logic_vector(15 downto 0);
    signal inc_2872 : std_logic_vector(15 downto 0);
    signal indvar_2702 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2931 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2919 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2723 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2913 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2716 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2893 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2906 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2709 : std_logic_vector(15 downto 0);
    signal mul59_2755 : std_logic_vector(15 downto 0);
    signal mul81_2777 : std_logic_vector(63 downto 0);
    signal mul83_2787 : std_logic_vector(63 downto 0);
    signal mul_2745 : std_logic_vector(15 downto 0);
    signal ptr_deref_2812_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2812_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2812_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2812_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2812_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2834_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2834_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2834_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2834_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2834_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2834_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_2626 : std_logic_vector(31 downto 0);
    signal shr135_2654 : std_logic_vector(15 downto 0);
    signal shr31136_2660 : std_logic_vector(15 downto 0);
    signal shr86_2798 : std_logic_vector(31 downto 0);
    signal shr90_2819 : std_logic_vector(63 downto 0);
    signal sub53_2750 : std_logic_vector(15 downto 0);
    signal sub66_2687 : std_logic_vector(15 downto 0);
    signal sub67_2760 : std_logic_vector(15 downto 0);
    signal sub_2676 : std_logic_vector(15 downto 0);
    signal tmp1_2735 : std_logic_vector(31 downto 0);
    signal tmp88_2813 : std_logic_vector(63 downto 0);
    signal type_cast_2624_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2652_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2658_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2669_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2680_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2706_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2708_wire : std_logic_vector(31 downto 0);
    signal type_cast_2713_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2715_wire : std_logic_vector(15 downto 0);
    signal type_cast_2720_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2722_wire : std_logic_vector(15 downto 0);
    signal type_cast_2726_wire : std_logic_vector(15 downto 0);
    signal type_cast_2728_wire : std_logic_vector(15 downto 0);
    signal type_cast_2733_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2796_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2817_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2823_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2844_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2862_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2870_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2890_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2909_wire : std_logic_vector(15 downto 0);
    signal type_cast_2912_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2916_wire : std_logic_vector(15 downto 0);
    signal type_cast_2918_wire : std_logic_vector(15 downto 0);
    signal type_cast_2922_wire : std_logic_vector(15 downto 0);
    signal type_cast_2924_wire : std_logic_vector(15 downto 0);
    signal type_cast_2929_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2937_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2807_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2807_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2807_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2807_resized_base_address <= "00000000000000";
    array_obj_ref_2830_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2830_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2830_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2830_resized_base_address <= "00000000000000";
    ptr_deref_2812_word_offset_0 <= "00000000000000";
    ptr_deref_2834_word_offset_0 <= "00000000000000";
    type_cast_2624_wire_constant <= "00000000000000000000000000010000";
    type_cast_2652_wire_constant <= "0000000000000010";
    type_cast_2658_wire_constant <= "0000000000000001";
    type_cast_2669_wire_constant <= "1111111111111111";
    type_cast_2680_wire_constant <= "1111111111111111";
    type_cast_2706_wire_constant <= "00000000000000000000000000000000";
    type_cast_2713_wire_constant <= "0000000000000000";
    type_cast_2720_wire_constant <= "0000000000000000";
    type_cast_2733_wire_constant <= "00000000000000000000000000000100";
    type_cast_2796_wire_constant <= "00000000000000000000000000000010";
    type_cast_2817_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_2823_wire_constant <= "0000000000000000000000000000000000111111111111111111111111111111";
    type_cast_2844_wire_constant <= "00000000000000000000000000000100";
    type_cast_2862_wire_constant <= "0000000000000100";
    type_cast_2870_wire_constant <= "0000000000000001";
    type_cast_2890_wire_constant <= "0000000000000000";
    type_cast_2912_wire_constant <= "0000000000000000";
    type_cast_2929_wire_constant <= "00000000000000000000000000000001";
    type_cast_2937_wire_constant <= "0000000000000001";
    phi_stmt_2702: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2706_wire_constant & type_cast_2708_wire;
      req <= phi_stmt_2702_req_0 & phi_stmt_2702_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2702",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2702_ack_0,
          idata => idata,
          odata => indvar_2702,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2702
    phi_stmt_2709: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2713_wire_constant & type_cast_2715_wire;
      req <= phi_stmt_2709_req_0 & phi_stmt_2709_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2709",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2709_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2709,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2709
    phi_stmt_2716: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2720_wire_constant & type_cast_2722_wire;
      req <= phi_stmt_2716_req_0 & phi_stmt_2716_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2716",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2716_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2716,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2716
    phi_stmt_2723: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2726_wire & type_cast_2728_wire;
      req <= phi_stmt_2723_req_0 & phi_stmt_2723_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2723",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2723_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2723,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2723
    phi_stmt_2906: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2909_wire & type_cast_2912_wire_constant;
      req <= phi_stmt_2906_req_0 & phi_stmt_2906_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2906",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2906_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2906,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2906
    phi_stmt_2913: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2916_wire & type_cast_2918_wire;
      req <= phi_stmt_2913_req_0 & phi_stmt_2913_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2913",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2913_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2913,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2913
    phi_stmt_2919: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2922_wire & type_cast_2924_wire;
      req <= phi_stmt_2919_req_0 & phi_stmt_2919_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2919",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2919_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2919,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2919
    -- flow-through select operator MUX_2892_inst
    input_dim1x_x2_2893 <= type_cast_2890_wire_constant when (cmp111_2877(0) /=  '0') else inc_2872;
    addr_of_2808_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2808_final_reg_req_0;
      addr_of_2808_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2808_final_reg_req_1;
      addr_of_2808_final_reg_ack_1<= rack(0);
      addr_of_2808_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2808_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2807_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx87_2809,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2831_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2831_final_reg_req_0;
      addr_of_2831_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2831_final_reg_req_1;
      addr_of_2831_final_reg_ack_1<= rack(0);
      addr_of_2831_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2831_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2830_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx92_2832,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2619_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2619_inst_req_0;
      type_cast_2619_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2619_inst_req_1;
      type_cast_2619_inst_ack_1<= rack(0);
      type_cast_2619_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2619_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_2616,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2620,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2632_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2632_inst_req_0;
      type_cast_2632_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2632_inst_req_1;
      type_cast_2632_inst_ack_1<= rack(0);
      type_cast_2632_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2632_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_2629,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_2633,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2690_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2690_inst_req_0;
      type_cast_2690_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2690_inst_req_1;
      type_cast_2690_inst_ack_1<= rack(0);
      type_cast_2690_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2690_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call22_2647,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_2691,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2694_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2694_inst_req_0;
      type_cast_2694_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2694_inst_req_1;
      type_cast_2694_inst_ack_1<= rack(0);
      type_cast_2694_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2694_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call20_2644,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv78_2695,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2698_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2698_inst_req_0;
      type_cast_2698_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2698_inst_req_1;
      type_cast_2698_inst_ack_1<= rack(0);
      type_cast_2698_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2698_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_2595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv99_2699,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2708_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2708_inst_req_0;
      type_cast_2708_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2708_inst_req_1;
      type_cast_2708_inst_ack_1<= rack(0);
      type_cast_2708_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2708_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2931,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2708_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2715_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2715_inst_req_0;
      type_cast_2715_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2715_inst_req_1;
      type_cast_2715_inst_ack_1<= rack(0);
      type_cast_2715_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2715_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2906,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2715_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2722_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2722_inst_req_0;
      type_cast_2722_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2722_inst_req_1;
      type_cast_2722_inst_ack_1<= rack(0);
      type_cast_2722_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2722_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2913,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2722_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2726_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2726_inst_req_0;
      type_cast_2726_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2726_inst_req_1;
      type_cast_2726_inst_ack_1<= rack(0);
      type_cast_2726_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2726_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add32_2665,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2726_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2728_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2728_inst_req_0;
      type_cast_2728_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2728_inst_req_1;
      type_cast_2728_inst_ack_1<= rack(0);
      type_cast_2728_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2728_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2919,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2728_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2763_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2763_inst_req_0;
      type_cast_2763_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2763_inst_req_1;
      type_cast_2763_inst_ack_1<= rack(0);
      type_cast_2763_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2763_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2709,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_2764,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2767_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2767_inst_req_0;
      type_cast_2767_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2767_inst_req_1;
      type_cast_2767_inst_ack_1<= rack(0);
      type_cast_2767_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2767_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub67_2760,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2768,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2771_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2771_inst_req_0;
      type_cast_2771_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2771_inst_req_1;
      type_cast_2771_inst_ack_1<= rack(0);
      type_cast_2771_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2771_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub53_2750,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_2772,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2801_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2801_inst_req_0;
      type_cast_2801_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2801_inst_req_1;
      type_cast_2801_inst_ack_1<= rack(0);
      type_cast_2801_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2801_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr86_2798,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2802,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2839_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2839_inst_req_0;
      type_cast_2839_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2839_inst_req_1;
      type_cast_2839_inst_ack_1<= rack(0);
      type_cast_2839_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2839_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2709,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_2840,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2880_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2880_inst_req_0;
      type_cast_2880_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2880_inst_req_1;
      type_cast_2880_inst_ack_1<= rack(0);
      type_cast_2880_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2880_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp111_2877,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc115_2881,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2909_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2909_inst_req_0;
      type_cast_2909_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2909_inst_req_1;
      type_cast_2909_inst_ack_1<= rack(0);
      type_cast_2909_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2909_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add103_2864,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2909_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2916_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2916_inst_req_0;
      type_cast_2916_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2916_inst_req_1;
      type_cast_2916_inst_ack_1<= rack(0);
      type_cast_2916_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2916_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2716,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2916_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2918_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2918_inst_req_0;
      type_cast_2918_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2918_inst_req_1;
      type_cast_2918_inst_ack_1<= rack(0);
      type_cast_2918_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2918_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2893,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2918_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2922_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2922_inst_req_0;
      type_cast_2922_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2922_inst_req_1;
      type_cast_2922_inst_ack_1<= rack(0);
      type_cast_2922_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2922_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2723,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2922_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2924_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2924_inst_req_0;
      type_cast_2924_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2924_inst_req_1;
      type_cast_2924_inst_ack_1<= rack(0);
      type_cast_2924_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2924_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc115x_xinput_dim0x_x2_2886,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2924_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2807_index_1_rename
    process(R_idxprom_2806_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2806_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2806_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2807_index_1_resize
    process(idxprom_2802) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2802;
      ov := iv(13 downto 0);
      R_idxprom_2806_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2807_root_address_inst
    process(array_obj_ref_2807_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2807_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2807_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2830_index_1_rename
    process(R_idxprom91_2829_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom91_2829_resized;
      ov(13 downto 0) := iv;
      R_idxprom91_2829_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2830_index_1_resize
    process(idxprom91_2825) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom91_2825;
      ov := iv(13 downto 0);
      R_idxprom91_2829_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2830_root_address_inst
    process(array_obj_ref_2830_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2830_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2830_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2812_addr_0
    process(ptr_deref_2812_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2812_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2812_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2812_base_resize
    process(arrayidx87_2809) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx87_2809;
      ov := iv(13 downto 0);
      ptr_deref_2812_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2812_gather_scatter
    process(ptr_deref_2812_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2812_data_0;
      ov(63 downto 0) := iv;
      tmp88_2813 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2812_root_address_inst
    process(ptr_deref_2812_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2812_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2812_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2834_addr_0
    process(ptr_deref_2834_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2834_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2834_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2834_base_resize
    process(arrayidx92_2832) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx92_2832;
      ov := iv(13 downto 0);
      ptr_deref_2834_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2834_gather_scatter
    process(tmp88_2813) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp88_2813;
      ov(63 downto 0) := iv;
      ptr_deref_2834_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2834_root_address_inst
    process(ptr_deref_2834_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2834_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2834_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2852_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2851;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2852_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2852_branch_req_0,
          ack0 => if_stmt_2852_branch_ack_0,
          ack1 => if_stmt_2852_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2899_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp121_2898;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2899_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2899_branch_req_0,
          ack0 => if_stmt_2899_branch_ack_0,
          ack1 => if_stmt_2899_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2664_inst
    process(shr135_2654, shr31136_2660) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr135_2654, shr31136_2660, tmp_var);
      add32_2665 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2670_inst
    process(call7_2601) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call7_2601, type_cast_2669_wire_constant, tmp_var);
      add50_2671 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2681_inst
    process(call9_2604) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call9_2604, type_cast_2680_wire_constant, tmp_var);
      add63_2682 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2749_inst
    process(sub_2676, mul_2745) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2676, mul_2745, tmp_var);
      sub53_2750 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2759_inst
    process(sub66_2687, mul59_2755) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub66_2687, mul59_2755, tmp_var);
      sub67_2760 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2863_inst
    process(input_dim2x_x1_2709) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2709, type_cast_2862_wire_constant, tmp_var);
      add103_2864 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2871_inst
    process(input_dim1x_x1_2716) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2716, type_cast_2870_wire_constant, tmp_var);
      inc_2872 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2885_inst
    process(inc115_2881, input_dim0x_x2_2723) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc115_2881, input_dim0x_x2_2723, tmp_var);
      inc115x_xinput_dim0x_x2_2886 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2739_inst
    process(add_2638, tmp1_2735) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_2638, tmp1_2735, tmp_var);
      add_src_0x_x0_2740 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2845_inst
    process(conv95_2840) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv95_2840, type_cast_2844_wire_constant, tmp_var);
      add96_2846 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2930_inst
    process(indvar_2702) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2702, type_cast_2929_wire_constant, tmp_var);
      indvarx_xnext_2931 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2781_inst
    process(mul81_2777, conv75_2768) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul81_2777, conv75_2768, tmp_var);
      add82_2782 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_2791_inst
    process(mul83_2787, conv70_2764) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul83_2787, conv70_2764, tmp_var);
      add84_2792 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_2824_inst
    process(shr90_2819) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr90_2819, type_cast_2823_wire_constant, tmp_var);
      idxprom91_2825 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2876_inst
    process(inc_2872, call1_2592) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_2872, call1_2592, tmp_var);
      cmp111_2877 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2897_inst
    process(inc115x_xinput_dim0x_x2_2886, call_2589) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc115x_xinput_dim0x_x2_2886, call_2589, tmp_var);
      cmp121_2898 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2653_inst
    process(call_2589) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2589, type_cast_2652_wire_constant, tmp_var);
      shr135_2654 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_2659_inst
    process(call_2589) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2589, type_cast_2658_wire_constant, tmp_var);
      shr31136_2660 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2797_inst
    process(add_src_0x_x0_2740) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2740, type_cast_2796_wire_constant, tmp_var);
      shr86_2798 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_2818_inst
    process(add84_2792) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add84_2792, type_cast_2817_wire_constant, tmp_var);
      shr90_2819 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2744_inst
    process(input_dim0x_x2_2723, call13_2610) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim0x_x2_2723, call13_2610, tmp_var);
      mul_2745 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2754_inst
    process(input_dim1x_x1_2716, call13_2610) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(input_dim1x_x1_2716, call13_2610, tmp_var);
      mul59_2755 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2734_inst
    process(indvar_2702) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2702, type_cast_2733_wire_constant, tmp_var);
      tmp1_2735 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2776_inst
    process(conv80_2772, conv78_2695) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv80_2772, conv78_2695, tmp_var);
      mul81_2777 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_2786_inst
    process(add82_2782, conv73_2691) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add82_2782, conv73_2691, tmp_var);
      mul83_2787 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_2637_inst
    process(shl_2626, conv17_2633) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_2626, conv17_2633, tmp_var);
      add_2638 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2625_inst
    process(conv_2620) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_2620, type_cast_2624_wire_constant, tmp_var);
      shl_2626 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2675_inst
    process(add50_2671, call14_2613) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add50_2671, call14_2613, tmp_var);
      sub_2676 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_2686_inst
    process(add63_2682, call14_2613) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(add63_2682, call14_2613, tmp_var);
      sub66_2687 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2850_inst
    process(add96_2846, conv99_2699) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add96_2846, conv99_2699, tmp_var);
      cmp_2851 <= tmp_var; --
    end process;
    -- shared split operator group (30) : array_obj_ref_2807_index_offset 
    ApIntAdd_group_30: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2806_scaled;
      array_obj_ref_2807_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2807_index_offset_req_0;
      array_obj_ref_2807_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2807_index_offset_req_1;
      array_obj_ref_2807_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_30_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : array_obj_ref_2830_index_offset 
    ApIntAdd_group_31: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom91_2829_scaled;
      array_obj_ref_2830_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2830_index_offset_req_0;
      array_obj_ref_2830_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2830_index_offset_req_1;
      array_obj_ref_2830_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_31_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared load operator group (0) : ptr_deref_2812_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2812_load_0_req_0;
      ptr_deref_2812_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2812_load_0_req_1;
      ptr_deref_2812_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2812_word_address_0;
      ptr_deref_2812_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2834_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2834_store_0_req_0;
      ptr_deref_2834_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2834_store_0_req_1;
      ptr_deref_2834_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2834_word_address_0;
      data_in <= ptr_deref_2834_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2588_inst RPIPE_Block3_start_2591_inst RPIPE_Block3_start_2594_inst RPIPE_Block3_start_2597_inst RPIPE_Block3_start_2600_inst RPIPE_Block3_start_2603_inst RPIPE_Block3_start_2606_inst RPIPE_Block3_start_2609_inst RPIPE_Block3_start_2612_inst RPIPE_Block3_start_2615_inst RPIPE_Block3_start_2628_inst RPIPE_Block3_start_2640_inst RPIPE_Block3_start_2643_inst RPIPE_Block3_start_2646_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 13 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 13 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 13 downto 0);
      signal guard_vector : std_logic_vector( 13 downto 0);
      constant outBUFs : IntegerArray(13 downto 0) := (13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(13 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false);
      constant guardBuffering: IntegerArray(13 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2);
      -- 
    begin -- 
      reqL_unguarded(13) <= RPIPE_Block3_start_2588_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Block3_start_2591_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block3_start_2594_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block3_start_2597_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block3_start_2600_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block3_start_2603_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block3_start_2606_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block3_start_2609_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block3_start_2612_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block3_start_2615_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block3_start_2628_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block3_start_2640_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block3_start_2643_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block3_start_2646_inst_req_0;
      RPIPE_Block3_start_2588_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Block3_start_2591_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block3_start_2594_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block3_start_2597_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block3_start_2600_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block3_start_2603_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block3_start_2606_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block3_start_2609_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block3_start_2612_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block3_start_2615_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block3_start_2628_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block3_start_2640_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block3_start_2643_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block3_start_2646_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(13) <= RPIPE_Block3_start_2588_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Block3_start_2591_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block3_start_2594_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block3_start_2597_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block3_start_2600_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block3_start_2603_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block3_start_2606_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block3_start_2609_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block3_start_2612_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block3_start_2615_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block3_start_2628_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block3_start_2640_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block3_start_2643_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block3_start_2646_inst_req_1;
      RPIPE_Block3_start_2588_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Block3_start_2591_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block3_start_2594_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block3_start_2597_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block3_start_2600_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block3_start_2603_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block3_start_2606_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block3_start_2609_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block3_start_2612_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block3_start_2615_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block3_start_2628_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block3_start_2640_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block3_start_2643_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block3_start_2646_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      call_2589 <= data_out(223 downto 208);
      call1_2592 <= data_out(207 downto 192);
      call3_2595 <= data_out(191 downto 176);
      call5_2598 <= data_out(175 downto 160);
      call7_2601 <= data_out(159 downto 144);
      call9_2604 <= data_out(143 downto 128);
      call11_2607 <= data_out(127 downto 112);
      call13_2610 <= data_out(111 downto 96);
      call14_2613 <= data_out(95 downto 80);
      call15_2616 <= data_out(79 downto 64);
      call16_2629 <= data_out(63 downto 48);
      call18_2641 <= data_out(47 downto 32);
      call20_2644 <= data_out(31 downto 16);
      call22_2647 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 14, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 14,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_2935_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_2935_inst_req_0;
      WPIPE_Block3_done_2935_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_2935_inst_req_1;
      WPIPE_Block3_done_2935_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2937_wire_constant;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_timer_resp_34_inst_req_0 : boolean;
  signal RPIPE_timer_resp_34_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_34_inst_req_1 : boolean;
  signal RPIPE_timer_resp_34_inst_ack_1 : boolean;
  signal WPIPE_timer_req_29_inst_req_0 : boolean;
  signal WPIPE_timer_req_29_inst_ack_0 : boolean;
  signal WPIPE_timer_req_29_inst_req_1 : boolean;
  signal WPIPE_timer_req_29_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_sample_start_
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Sample/rr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/$entry
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_sample_start_
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Sample/req
      -- 
    req_13_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_13_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => WPIPE_timer_req_29_inst_req_0); -- 
    rr_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => RPIPE_timer_resp_34_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_sample_completed_
      -- CP-element group 1: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_update_start_
      -- CP-element group 1: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Sample/ack
      -- CP-element group 1: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Update/$entry
      -- CP-element group 1: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Update/req
      -- 
    ack_14_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_29_inst_ack_0, ack => timer_CP_0_elements(1)); -- 
    req_18_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_18_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(1), ack => WPIPE_timer_req_29_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_update_completed_
      -- CP-element group 2: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Update/$exit
      -- CP-element group 2: 	 assign_stmt_32_to_assign_stmt_35/WPIPE_timer_req_29_Update/ack
      -- 
    ack_19_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_29_inst_ack_1, ack => timer_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_sample_completed_
      -- CP-element group 3: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_update_start_
      -- CP-element group 3: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Sample/ra
      -- CP-element group 3: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Update/$entry
      -- CP-element group 3: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Update/cr
      -- 
    ra_28_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_34_inst_ack_0, ack => timer_CP_0_elements(3)); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(3), ack => RPIPE_timer_resp_34_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_update_completed_
      -- CP-element group 4: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Update/$exit
      -- CP-element group 4: 	 assign_stmt_32_to_assign_stmt_35/RPIPE_timer_resp_34_Update/ca
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_34_inst_ack_1, ack => timer_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_32_to_assign_stmt_35/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_0_elements(2) & timer_CP_0_elements(4);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_31_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_31_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_34_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_34_inst_req_0;
      RPIPE_timer_resp_34_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_34_inst_req_1;
      RPIPE_timer_resp_34_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_29_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_29_inst_req_0;
      WPIPE_timer_req_29_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_29_inst_req_1;
      WPIPE_timer_req_29_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_31_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    timer_req_pipe_read_data: out std_logic_vector(0 downto 0);
    timer_req_pipe_read_req : in std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : out std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data: in std_logic_vector(63 downto 0);
    timer_resp_pipe_write_req : in std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(4 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(18 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(10 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(0 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(4 downto 4),
      memory_space_2_sr_ack => memory_space_2_sr_ack(4 downto 4),
      memory_space_2_sr_addr => memory_space_2_sr_addr(69 downto 56),
      memory_space_2_sr_data => memory_space_2_sr_data(319 downto 256),
      memory_space_2_sr_tag => memory_space_2_sr_tag(94 downto 76),
      memory_space_2_sc_req => memory_space_2_sc_req(4 downto 4),
      memory_space_2_sc_ack => memory_space_2_sc_ack(4 downto 4),
      memory_space_2_sc_tag => memory_space_2_sc_tag(4 downto 4),
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(3 downto 3),
      memory_space_0_lr_ack => memory_space_0_lr_ack(3 downto 3),
      memory_space_0_lr_addr => memory_space_0_lr_addr(55 downto 42),
      memory_space_0_lr_tag => memory_space_0_lr_tag(75 downto 57),
      memory_space_0_lc_req => memory_space_0_lc_req(3 downto 3),
      memory_space_0_lc_ack => memory_space_0_lc_ack(3 downto 3),
      memory_space_0_lc_data => memory_space_0_lc_data(255 downto 192),
      memory_space_0_lc_tag => memory_space_0_lc_tag(3 downto 3),
      memory_space_2_sr_req => memory_space_2_sr_req(3 downto 3),
      memory_space_2_sr_ack => memory_space_2_sr_ack(3 downto 3),
      memory_space_2_sr_addr => memory_space_2_sr_addr(55 downto 42),
      memory_space_2_sr_data => memory_space_2_sr_data(255 downto 192),
      memory_space_2_sr_tag => memory_space_2_sr_tag(75 downto 57),
      memory_space_2_sc_req => memory_space_2_sc_req(3 downto 3),
      memory_space_2_sc_ack => memory_space_2_sc_ack(3 downto 3),
      memory_space_2_sc_tag => memory_space_2_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(2 downto 2),
      memory_space_0_lr_ack => memory_space_0_lr_ack(2 downto 2),
      memory_space_0_lr_addr => memory_space_0_lr_addr(41 downto 28),
      memory_space_0_lr_tag => memory_space_0_lr_tag(56 downto 38),
      memory_space_0_lc_req => memory_space_0_lc_req(2 downto 2),
      memory_space_0_lc_ack => memory_space_0_lc_ack(2 downto 2),
      memory_space_0_lc_data => memory_space_0_lc_data(191 downto 128),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 2),
      memory_space_2_sr_req => memory_space_2_sr_req(2 downto 2),
      memory_space_2_sr_ack => memory_space_2_sr_ack(2 downto 2),
      memory_space_2_sr_addr => memory_space_2_sr_addr(41 downto 28),
      memory_space_2_sr_data => memory_space_2_sr_data(191 downto 128),
      memory_space_2_sr_tag => memory_space_2_sr_tag(56 downto 38),
      memory_space_2_sc_req => memory_space_2_sc_req(2 downto 2),
      memory_space_2_sc_ack => memory_space_2_sc_ack(2 downto 2),
      memory_space_2_sc_tag => memory_space_2_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(27 downto 14),
      memory_space_0_lr_tag => memory_space_0_lr_tag(37 downto 19),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(127 downto 64),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 1),
      memory_space_2_sr_req => memory_space_2_sr_req(1 downto 1),
      memory_space_2_sr_ack => memory_space_2_sr_ack(1 downto 1),
      memory_space_2_sr_addr => memory_space_2_sr_addr(27 downto 14),
      memory_space_2_sr_data => memory_space_2_sr_data(127 downto 64),
      memory_space_2_sr_tag => memory_space_2_sr_tag(37 downto 19),
      memory_space_2_sc_req => memory_space_2_sc_req(1 downto 1),
      memory_space_2_sc_ack => memory_space_2_sc_ack(1 downto 1),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 1),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(13 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(18 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_1: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
