-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_26_start: Boolean;
  signal timer_CP_26_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_20_load_0_req_0 : boolean;
  signal LOAD_count_20_load_0_ack_0 : boolean;
  signal LOAD_count_20_load_0_req_1 : boolean;
  signal LOAD_count_20_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_26_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_26_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_26_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_26_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_26: Block -- control-path 
    signal timer_CP_26_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_26_elements(0) <= timer_CP_26_start;
    timer_CP_26_symbol <= timer_CP_26_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_21/$entry
      -- CP-element group 0: 	 assign_stmt_21/LOAD_count_20_sample_start_
      -- CP-element group 0: 	 assign_stmt_21/LOAD_count_20_update_start_
      -- CP-element group 0: 	 assign_stmt_21/LOAD_count_20_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_21/LOAD_count_20_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_21/LOAD_count_20_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_21/LOAD_count_20_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_21/LOAD_count_20_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_21/LOAD_count_20_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_21/LOAD_count_20_Update/$entry
      -- CP-element group 0: 	 assign_stmt_21/LOAD_count_20_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_21/LOAD_count_20_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_21/LOAD_count_20_Update/word_access_complete/word_0/cr
      -- 
    cr_58_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_58_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_26_elements(0), ack => LOAD_count_20_load_0_req_1); -- 
    rr_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_26_elements(0), ack => LOAD_count_20_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_21/LOAD_count_20_sample_completed_
      -- CP-element group 1: 	 assign_stmt_21/LOAD_count_20_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_21/LOAD_count_20_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_21/LOAD_count_20_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_21/LOAD_count_20_Sample/word_access_start/word_0/ra
      -- 
    ra_48_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_20_load_0_ack_0, ack => timer_CP_26_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_21/$exit
      -- CP-element group 2: 	 assign_stmt_21/LOAD_count_20_update_completed_
      -- CP-element group 2: 	 assign_stmt_21/LOAD_count_20_Update/$exit
      -- CP-element group 2: 	 assign_stmt_21/LOAD_count_20_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_21/LOAD_count_20_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_21/LOAD_count_20_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_21/LOAD_count_20_Update/LOAD_count_20_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_21/LOAD_count_20_Update/LOAD_count_20_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_21/LOAD_count_20_Update/LOAD_count_20_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_21/LOAD_count_20_Update/LOAD_count_20_Merge/merge_ack
      -- 
    ca_59_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_20_load_0_ack_1, ack => timer_CP_26_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_20_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_20_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_20_word_address_0 <= "0";
    -- equivalence LOAD_count_20_gather_scatter
    process(LOAD_count_20_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_20_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_20_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_20_load_0_req_0;
      LOAD_count_20_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_20_load_0_req_1;
      LOAD_count_20_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_20_word_address_0;
      LOAD_count_20_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(0 downto 0),
          mtag => memory_space_1_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_65_start: Boolean;
  signal timerDaemon_CP_65_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_25_branch_req_0 : boolean;
  signal phi_stmt_27_req_1 : boolean;
  signal phi_stmt_27_req_0 : boolean;
  signal phi_stmt_27_ack_0 : boolean;
  signal ADD_u64_u64_33_inst_req_0 : boolean;
  signal ADD_u64_u64_33_inst_ack_0 : boolean;
  signal ADD_u64_u64_33_inst_req_1 : boolean;
  signal ADD_u64_u64_33_inst_ack_1 : boolean;
  signal STORE_count_35_store_0_req_0 : boolean;
  signal STORE_count_35_store_0_ack_0 : boolean;
  signal STORE_count_35_store_0_req_1 : boolean;
  signal STORE_count_35_store_0_ack_1 : boolean;
  signal do_while_stmt_25_branch_ack_0 : boolean;
  signal do_while_stmt_25_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_65_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_65_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_65_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_65_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_65: Block -- control-path 
    signal timerDaemon_CP_65_elements: BooleanArray(39 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_65_elements(0) <= timerDaemon_CP_65_start;
    timerDaemon_CP_65_symbol <= timerDaemon_CP_65_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_24/$entry
      -- CP-element group 0: 	 branch_block_stmt_24/branch_block_stmt_24__entry__
      -- CP-element group 0: 	 branch_block_stmt_24/do_while_stmt_25__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	39 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_24/$exit
      -- CP-element group 1: 	 branch_block_stmt_24/branch_block_stmt_24__exit__
      -- CP-element group 1: 	 branch_block_stmt_24/do_while_stmt_25__exit__
      -- 
    timerDaemon_CP_65_elements(1) <= timerDaemon_CP_65_elements(39);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_24/do_while_stmt_25/$entry
      -- CP-element group 2: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25__entry__
      -- 
    timerDaemon_CP_65_elements(2) <= timerDaemon_CP_65_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	39 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25__exit__
      -- 
    -- Element group timerDaemon_CP_65_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_24/do_while_stmt_25/loop_back
      -- 
    -- Element group timerDaemon_CP_65_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	37 
    -- CP-element group 5: 	38 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_24/do_while_stmt_25/condition_done
      -- CP-element group 5: 	 branch_block_stmt_24/do_while_stmt_25/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_24/do_while_stmt_25/loop_taken/$entry
      -- 
    timerDaemon_CP_65_elements(5) <= timerDaemon_CP_65_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	36 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_24/do_while_stmt_25/loop_body_done
      -- 
    timerDaemon_CP_65_elements(6) <= timerDaemon_CP_65_elements(36);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_65_elements(7) <= timerDaemon_CP_65_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_65_elements(8) <= timerDaemon_CP_65_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	31 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	35 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_root_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/loop_body_start
      -- 
    -- Element group timerDaemon_CP_65_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	35 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/condition_evaluated
      -- 
    condition_evaluated_89_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_89_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_65_elements(10), ack => do_while_stmt_25_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_65_elements(15) & timerDaemon_CP_65_elements(35);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_65_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/phi_stmt_27_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_65_elements(12) & timerDaemon_CP_65_elements(15);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_65_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/phi_stmt_27_sample_start_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_65_elements(9) & timerDaemon_CP_65_elements(14);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_65_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	33 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/phi_stmt_27_update_start_
      -- CP-element group 13: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/phi_stmt_27_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_65_elements(9) & timerDaemon_CP_65_elements(33);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_65_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/phi_stmt_27_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/phi_stmt_27_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_65_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	31 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/phi_stmt_27_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/phi_stmt_27_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_65_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/phi_stmt_27_loopback_trigger
      -- 
    timerDaemon_CP_65_elements(16) <= timerDaemon_CP_65_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/phi_stmt_27_loopback_sample_req
      -- CP-element group 17: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/phi_stmt_27_loopback_sample_req_ps
      -- 
    phi_stmt_27_loopback_sample_req_104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_27_loopback_sample_req_104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_65_elements(17), ack => phi_stmt_27_req_1); -- 
    -- Element group timerDaemon_CP_65_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/phi_stmt_27_entry_trigger
      -- 
    timerDaemon_CP_65_elements(18) <= timerDaemon_CP_65_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/phi_stmt_27_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/phi_stmt_27_entry_sample_req_ps
      -- 
    phi_stmt_27_entry_sample_req_107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_27_entry_sample_req_107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_65_elements(19), ack => phi_stmt_27_req_0); -- 
    -- Element group timerDaemon_CP_65_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/phi_stmt_27_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/phi_stmt_27_phi_mux_ack_ps
      -- 
    phi_stmt_27_phi_mux_ack_110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_27_ack_0, ack => timerDaemon_CP_65_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/type_cast_30_sample_start__ps
      -- CP-element group 21: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/type_cast_30_sample_completed__ps
      -- CP-element group 21: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/type_cast_30_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/type_cast_30_sample_completed_
      -- 
    -- Element group timerDaemon_CP_65_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/type_cast_30_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/type_cast_30_update_start_
      -- 
    -- Element group timerDaemon_CP_65_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/type_cast_30_update_completed__ps
      -- 
    timerDaemon_CP_65_elements(23) <= timerDaemon_CP_65_elements(24);
    -- CP-element group 24:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	23 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/type_cast_30_update_completed_
      -- 
    -- Element group timerDaemon_CP_65_elements(24) is a control-delay.
    cp_element_24_delay: control_delay_element  generic map(name => " 24_delay", delay_value => 1)  port map(req => timerDaemon_CP_65_elements(22), ack => timerDaemon_CP_65_elements(24), clk => clk, reset =>reset);
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/ADD_u64_u64_33_sample_start__ps
      -- 
    -- Element group timerDaemon_CP_65_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/ADD_u64_u64_33_update_start__ps
      -- 
    -- Element group timerDaemon_CP_65_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/ADD_u64_u64_33_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/ADD_u64_u64_33_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/ADD_u64_u64_33_Sample/rr
      -- 
    rr_131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_65_elements(27), ack => ADD_u64_u64_33_inst_req_0); -- 
    timerDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_65_elements(25) & timerDaemon_CP_65_elements(29);
      gj_timerDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_65_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/ADD_u64_u64_33_update_start_
      -- CP-element group 28: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/ADD_u64_u64_33_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/ADD_u64_u64_33_Update/cr
      -- 
    cr_136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_65_elements(28), ack => ADD_u64_u64_33_inst_req_1); -- 
    timerDaemon_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_65_elements(26) & timerDaemon_CP_65_elements(30);
      gj_timerDaemon_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_65_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/ADD_u64_u64_33_sample_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/ADD_u64_u64_33_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/ADD_u64_u64_33_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/ADD_u64_u64_33_Sample/ra
      -- 
    ra_132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_33_inst_ack_0, ack => timerDaemon_CP_65_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/ADD_u64_u64_33_update_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/ADD_u64_u64_33_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/ADD_u64_u64_33_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/ADD_u64_u64_33_Update/ca
      -- 
    ca_137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_33_inst_ack_1, ack => timerDaemon_CP_65_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	9 
    -- CP-element group 31: 	15 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Sample/STORE_count_35_Split/$entry
      -- CP-element group 31: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Sample/STORE_count_35_Split/$exit
      -- CP-element group 31: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Sample/STORE_count_35_Split/split_req
      -- CP-element group 31: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Sample/STORE_count_35_Split/split_ack
      -- CP-element group 31: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Sample/word_access_start/word_0/rr
      -- 
    rr_159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_65_elements(31), ack => STORE_count_35_store_0_req_0); -- 
    timerDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 3,1 => 3,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_65_elements(9) & timerDaemon_CP_65_elements(15) & timerDaemon_CP_65_elements(33);
      gj_timerDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_65_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_update_start_
      -- CP-element group 32: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Update/word_access_complete/$entry
      -- CP-element group 32: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Update/word_access_complete/word_0/$entry
      -- CP-element group 32: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Update/word_access_complete/word_0/cr
      -- 
    cr_170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_65_elements(32), ack => STORE_count_35_store_0_req_1); -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= timerDaemon_CP_65_elements(34);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_65_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: 	13 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Sample/word_access_start/$exit
      -- CP-element group 33: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Sample/word_access_start/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Sample/word_access_start/word_0/ra
      -- 
    ra_160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_35_store_0_ack_0, ack => timerDaemon_CP_65_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Update/word_access_complete/$exit
      -- CP-element group 34: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Update/word_access_complete/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/STORE_count_35_Update/word_access_complete/word_0/ca
      -- 
    ca_171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_35_store_0_ack_1, ack => timerDaemon_CP_65_elements(34)); -- 
    -- CP-element group 35:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	10 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_65_elements(35) is a control-delay.
    cp_element_35_delay: control_delay_element  generic map(name => " 35_delay", delay_value => 1)  port map(req => timerDaemon_CP_65_elements(9), ack => timerDaemon_CP_65_elements(35), clk => clk, reset =>reset);
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	6 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_24/do_while_stmt_25/do_while_stmt_25_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_65_elements(14) & timerDaemon_CP_65_elements(34);
      gj_timerDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_65_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	5 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_24/do_while_stmt_25/loop_exit/$exit
      -- CP-element group 37: 	 branch_block_stmt_24/do_while_stmt_25/loop_exit/ack
      -- 
    ack_176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_25_branch_ack_0, ack => timerDaemon_CP_65_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	5 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_24/do_while_stmt_25/loop_taken/$exit
      -- CP-element group 38: 	 branch_block_stmt_24/do_while_stmt_25/loop_taken/ack
      -- 
    ack_180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_25_branch_ack_1, ack => timerDaemon_CP_65_elements(38)); -- 
    -- CP-element group 39:  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	3 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	1 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_24/do_while_stmt_25/$exit
      -- 
    timerDaemon_CP_65_elements(39) <= timerDaemon_CP_65_elements(3);
    timerDaemon_do_while_stmt_25_terminator_181: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_25_terminator_181", max_iterations_in_flight =>3) 
      port map(loop_body_exit => timerDaemon_CP_65_elements(6),loop_continue => timerDaemon_CP_65_elements(38),loop_terminate => timerDaemon_CP_65_elements(37),loop_back => timerDaemon_CP_65_elements(4),loop_exit => timerDaemon_CP_65_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_27_phi_seq_138_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_65_elements(18);
      timerDaemon_CP_65_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_65_elements(21);
      timerDaemon_CP_65_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_65_elements(23);
      timerDaemon_CP_65_elements(19) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_65_elements(16);
      timerDaemon_CP_65_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_65_elements(29);
      timerDaemon_CP_65_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_65_elements(30);
      timerDaemon_CP_65_elements(17) <= phi_mux_reqs(1);
      phi_stmt_27_phi_seq_138 : phi_sequencer_v2-- 
        generic map (place_capacity => 3, ntriggers => 2, name => "phi_stmt_27_phi_seq_138") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_65_elements(11), 
          phi_sample_ack => timerDaemon_CP_65_elements(14), 
          phi_update_req => timerDaemon_CP_65_elements(13), 
          phi_update_ack => timerDaemon_CP_65_elements(15), 
          phi_mux_ack => timerDaemon_CP_65_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_90_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_65_elements(7);
        preds(1)  <= timerDaemon_CP_65_elements(8);
        entry_tmerge_90 : transition_merge -- 
          generic map(name => " entry_tmerge_90")
          port map (preds => preds, symbol_out => timerDaemon_CP_65_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u64_u64_33_wire : std_logic_vector(63 downto 0);
    signal STORE_count_35_data_0 : std_logic_vector(63 downto 0);
    signal STORE_count_35_word_address_0 : std_logic_vector(0 downto 0);
    signal konst_32_wire_constant : std_logic_vector(63 downto 0);
    signal konst_39_wire_constant : std_logic_vector(0 downto 0);
    signal ncount_27 : std_logic_vector(63 downto 0);
    signal type_cast_30_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_count_35_word_address_0 <= "0";
    konst_32_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_39_wire_constant <= "1";
    type_cast_30_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_27: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_30_wire_constant & ADD_u64_u64_33_wire;
      req <= phi_stmt_27_req_0 & phi_stmt_27_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_27",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_27_ack_0,
          idata => idata,
          odata => ncount_27,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_27
    -- equivalence STORE_count_35_gather_scatter
    process(ncount_27) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ncount_27;
      ov(63 downto 0) := iv;
      STORE_count_35_data_0 <= ov(63 downto 0);
      --
    end process;
    do_while_stmt_25_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_39_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_25_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_25_branch_req_0,
          ack0 => do_while_stmt_25_branch_ack_0,
          ack1 => do_while_stmt_25_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u64_u64_33_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ncount_27;
      ADD_u64_u64_33_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_33_inst_req_0;
      ADD_u64_u64_33_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_33_inst_req_1;
      ADD_u64_u64_33_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared store operator group (0) : STORE_count_35_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_count_35_store_0_req_0;
      STORE_count_35_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_count_35_store_0_req_1;
      STORE_count_35_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_count_35_word_address_0;
      data_in <= STORE_count_35_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(0 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(14 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(14 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    Zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    Zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad;
architecture zeropad_arch of zeropad is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad_CP_182_start: Boolean;
  signal zeropad_CP_182_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal W_ifx_xthen191_exec_guard_829_delayed_1_0_865_inst_ack_0 : boolean;
  signal W_output_byte_countx_x0_1017_delayed_2_0_1150_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1430_inst_ack_1 : boolean;
  signal phi_stmt_610_req_1 : boolean;
  signal type_cast_871_inst_ack_0 : boolean;
  signal type_cast_603_inst_ack_0 : boolean;
  signal MUX_1131_inst_ack_0 : boolean;
  signal type_cast_603_inst_req_0 : boolean;
  signal type_cast_613_inst_req_0 : boolean;
  signal W_ifx_xthen191_exec_guard_823_delayed_1_0_856_inst_req_1 : boolean;
  signal array_obj_ref_789_index_offset_ack_1 : boolean;
  signal type_cast_871_inst_ack_1 : boolean;
  signal W_ifx_xthen191_exec_guard_850_delayed_1_0_897_inst_ack_0 : boolean;
  signal addr_of_790_final_reg_req_1 : boolean;
  signal ptr_deref_1192_store_0_ack_0 : boolean;
  signal W_ifx_xthen191_exec_guard_850_delayed_1_0_897_inst_req_1 : boolean;
  signal W_ifx_xthen191_exec_guard_850_delayed_1_0_897_inst_ack_1 : boolean;
  signal phi_stmt_590_ack_0 : boolean;
  signal target_out_offsetx_x1_at_entry_539_599_buf_ack_1 : boolean;
  signal target_out_offsetx_x1_at_entry_539_599_buf_req_1 : boolean;
  signal ptr_deref_1192_store_0_req_0 : boolean;
  signal array_obj_ref_789_index_offset_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_59_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_59_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_59_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_59_inst_ack_1 : boolean;
  signal ptr_deref_798_load_0_ack_1 : boolean;
  signal type_cast_915_inst_req_1 : boolean;
  signal type_cast_593_inst_ack_1 : boolean;
  signal phi_stmt_605_req_0 : boolean;
  signal target_out_offsetx_x1_at_entry_539_599_buf_ack_0 : boolean;
  signal ptr_deref_798_load_0_req_1 : boolean;
  signal W_ifx_xthen191_exec_guard_829_delayed_1_0_865_inst_req_1 : boolean;
  signal W_ifx_xthen191_exec_guard_850_delayed_1_0_897_inst_req_0 : boolean;
  signal type_cast_593_inst_req_1 : boolean;
  signal MUX_1113_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1445_inst_req_0 : boolean;
  signal type_cast_613_inst_req_1 : boolean;
  signal phi_stmt_610_req_0 : boolean;
  signal type_cast_613_inst_ack_0 : boolean;
  signal W_o1x_x1_860_delayed_1_0_909_inst_ack_0 : boolean;
  signal W_o1x_x1_860_delayed_1_0_909_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1605_inst_req_0 : boolean;
  signal type_cast_613_inst_ack_1 : boolean;
  signal phi_stmt_610_ack_0 : boolean;
  signal W_ifx_xthen191_exec_guard_829_delayed_1_0_865_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue208_exec_guard_863_delayed_1_0_917_inst_ack_1 : boolean;
  signal W_ifx_xthen191_exec_guard_823_delayed_1_0_856_inst_ack_1 : boolean;
  signal W_ifx_xthen191_exec_guard_829_delayed_1_0_865_inst_ack_1 : boolean;
  signal phi_stmt_595_req_0 : boolean;
  signal type_cast_593_inst_ack_0 : boolean;
  signal type_cast_593_inst_req_0 : boolean;
  signal phi_stmt_590_req_1 : boolean;
  signal ptr_deref_491_load_0_ack_0 : boolean;
  signal ptr_deref_491_load_0_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_45_inst_req_0 : boolean;
  signal type_cast_1091_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_45_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_45_inst_req_1 : boolean;
  signal type_cast_598_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_45_inst_ack_1 : boolean;
  signal target_out_offsetx_x1_at_entry_539_599_buf_req_0 : boolean;
  signal type_cast_50_inst_req_0 : boolean;
  signal type_cast_50_inst_ack_0 : boolean;
  signal type_cast_50_inst_req_1 : boolean;
  signal type_cast_598_inst_req_1 : boolean;
  signal type_cast_50_inst_ack_1 : boolean;
  signal addr_of_284_final_reg_req_0 : boolean;
  signal addr_of_284_final_reg_ack_0 : boolean;
  signal addr_of_284_final_reg_req_1 : boolean;
  signal addr_of_284_final_reg_ack_1 : boolean;
  signal type_cast_1091_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_287_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_287_inst_ack_0 : boolean;
  signal addr_of_790_final_reg_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_287_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_287_inst_ack_1 : boolean;
  signal type_cast_915_inst_req_0 : boolean;
  signal type_cast_63_inst_req_0 : boolean;
  signal type_cast_63_inst_ack_0 : boolean;
  signal phi_stmt_600_ack_0 : boolean;
  signal type_cast_63_inst_req_1 : boolean;
  signal type_cast_63_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_71_inst_req_0 : boolean;
  signal type_cast_598_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_71_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_71_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_71_inst_ack_1 : boolean;
  signal type_cast_75_inst_req_0 : boolean;
  signal type_cast_598_inst_req_0 : boolean;
  signal type_cast_75_inst_ack_0 : boolean;
  signal type_cast_75_inst_req_1 : boolean;
  signal type_cast_75_inst_ack_1 : boolean;
  signal type_cast_608_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_84_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_84_inst_ack_0 : boolean;
  signal type_cast_608_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_84_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_84_inst_ack_1 : boolean;
  signal phi_stmt_605_ack_0 : boolean;
  signal type_cast_915_inst_ack_1 : boolean;
  signal type_cast_88_inst_req_0 : boolean;
  signal type_cast_88_inst_ack_0 : boolean;
  signal type_cast_88_inst_req_1 : boolean;
  signal type_cast_88_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_96_inst_req_0 : boolean;
  signal type_cast_1210_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_96_inst_ack_0 : boolean;
  signal phi_stmt_590_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_96_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_96_inst_ack_1 : boolean;
  signal type_cast_100_inst_req_0 : boolean;
  signal type_cast_100_inst_ack_0 : boolean;
  signal type_cast_100_inst_req_1 : boolean;
  signal type_cast_100_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_109_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_109_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_109_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_109_inst_ack_1 : boolean;
  signal type_cast_113_inst_req_0 : boolean;
  signal type_cast_113_inst_ack_0 : boolean;
  signal type_cast_113_inst_req_1 : boolean;
  signal type_cast_113_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_121_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_121_inst_ack_0 : boolean;
  signal type_cast_608_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_121_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_121_inst_ack_1 : boolean;
  signal type_cast_126_inst_req_0 : boolean;
  signal type_cast_126_inst_ack_0 : boolean;
  signal type_cast_126_inst_req_1 : boolean;
  signal type_cast_126_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_135_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_135_inst_ack_0 : boolean;
  signal type_cast_608_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_135_inst_req_1 : boolean;
  signal MUX_1131_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_135_inst_ack_1 : boolean;
  signal array_obj_ref_1187_index_offset_ack_1 : boolean;
  signal W_ifx_xthen191_exec_guard_838_delayed_1_0_880_inst_req_0 : boolean;
  signal type_cast_139_inst_req_0 : boolean;
  signal type_cast_139_inst_ack_0 : boolean;
  signal type_cast_139_inst_req_1 : boolean;
  signal type_cast_139_inst_ack_1 : boolean;
  signal type_cast_871_inst_req_1 : boolean;
  signal array_obj_ref_789_index_offset_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_147_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_147_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_147_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_147_inst_ack_1 : boolean;
  signal W_ifx_xthen191_exec_guard_838_delayed_1_0_880_inst_ack_0 : boolean;
  signal phi_stmt_600_req_1 : boolean;
  signal type_cast_151_inst_req_0 : boolean;
  signal phi_stmt_595_ack_0 : boolean;
  signal type_cast_151_inst_ack_0 : boolean;
  signal type_cast_151_inst_req_1 : boolean;
  signal type_cast_151_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_160_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_160_inst_ack_0 : boolean;
  signal do_while_stmt_588_branch_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_160_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_160_inst_ack_1 : boolean;
  signal W_ifx_xthen191_exec_guard_838_delayed_1_0_880_inst_req_1 : boolean;
  signal type_cast_164_inst_req_0 : boolean;
  signal type_cast_164_inst_ack_0 : boolean;
  signal type_cast_164_inst_req_1 : boolean;
  signal type_cast_164_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_172_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_172_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_172_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_172_inst_ack_1 : boolean;
  signal type_cast_603_inst_ack_1 : boolean;
  signal W_ifx_xthen191_exec_guard_838_delayed_1_0_880_inst_ack_1 : boolean;
  signal type_cast_176_inst_req_0 : boolean;
  signal type_cast_176_inst_ack_0 : boolean;
  signal type_cast_176_inst_req_1 : boolean;
  signal type_cast_176_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_185_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_185_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_185_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_185_inst_ack_1 : boolean;
  signal type_cast_603_inst_req_1 : boolean;
  signal type_cast_189_inst_req_0 : boolean;
  signal type_cast_189_inst_ack_0 : boolean;
  signal type_cast_189_inst_req_1 : boolean;
  signal type_cast_189_inst_ack_1 : boolean;
  signal phi_stmt_595_req_1 : boolean;
  signal type_cast_208_inst_req_0 : boolean;
  signal type_cast_208_inst_ack_0 : boolean;
  signal type_cast_208_inst_req_1 : boolean;
  signal type_cast_208_inst_ack_1 : boolean;
  signal array_obj_ref_789_index_offset_req_1 : boolean;
  signal type_cast_212_inst_req_0 : boolean;
  signal type_cast_212_inst_ack_0 : boolean;
  signal phi_stmt_600_req_0 : boolean;
  signal type_cast_212_inst_req_1 : boolean;
  signal type_cast_212_inst_ack_1 : boolean;
  signal ptr_deref_491_load_0_ack_1 : boolean;
  signal phi_stmt_605_req_1 : boolean;
  signal type_cast_871_inst_req_0 : boolean;
  signal type_cast_1530_inst_req_1 : boolean;
  signal ptr_deref_491_load_0_req_1 : boolean;
  signal if_stmt_231_branch_req_0 : boolean;
  signal if_stmt_231_branch_ack_1 : boolean;
  signal if_stmt_231_branch_ack_0 : boolean;
  signal addr_of_790_final_reg_ack_1 : boolean;
  signal W_ifx_xthen180_exec_guard_768_delayed_6_0_792_inst_req_0 : boolean;
  signal array_obj_ref_283_index_offset_req_0 : boolean;
  signal array_obj_ref_283_index_offset_ack_0 : boolean;
  signal array_obj_ref_283_index_offset_req_1 : boolean;
  signal array_obj_ref_283_index_offset_ack_1 : boolean;
  signal type_cast_291_inst_req_0 : boolean;
  signal type_cast_291_inst_ack_0 : boolean;
  signal type_cast_291_inst_req_1 : boolean;
  signal type_cast_291_inst_ack_1 : boolean;
  signal MUX_1113_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_300_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_300_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_300_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_300_inst_ack_1 : boolean;
  signal W_ifx_xthen191_exec_guard_845_delayed_1_0_889_inst_req_0 : boolean;
  signal W_ifx_xthen191_exec_guard_845_delayed_1_0_889_inst_ack_0 : boolean;
  signal type_cast_304_inst_req_0 : boolean;
  signal type_cast_304_inst_ack_0 : boolean;
  signal type_cast_1530_inst_ack_1 : boolean;
  signal type_cast_304_inst_req_1 : boolean;
  signal type_cast_304_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_318_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_318_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_318_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_318_inst_ack_1 : boolean;
  signal W_ifx_xthen180_exec_guard_768_delayed_6_0_792_inst_ack_0 : boolean;
  signal W_ifx_xthen191_exec_guard_845_delayed_1_0_889_inst_req_1 : boolean;
  signal type_cast_322_inst_req_0 : boolean;
  signal type_cast_322_inst_ack_0 : boolean;
  signal type_cast_322_inst_req_1 : boolean;
  signal type_cast_322_inst_ack_1 : boolean;
  signal ptr_deref_798_load_0_req_0 : boolean;
  signal ptr_deref_798_load_0_ack_0 : boolean;
  signal W_ifx_xthen191_exec_guard_845_delayed_1_0_889_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_336_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_336_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_336_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_336_inst_ack_1 : boolean;
  signal type_cast_340_inst_req_0 : boolean;
  signal type_cast_340_inst_ack_0 : boolean;
  signal type_cast_340_inst_req_1 : boolean;
  signal type_cast_340_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_354_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_354_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_354_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_354_inst_ack_1 : boolean;
  signal type_cast_358_inst_req_0 : boolean;
  signal type_cast_358_inst_ack_0 : boolean;
  signal type_cast_358_inst_req_1 : boolean;
  signal type_cast_358_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_372_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_372_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_372_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_372_inst_ack_1 : boolean;
  signal type_cast_376_inst_req_0 : boolean;
  signal type_cast_376_inst_ack_0 : boolean;
  signal type_cast_376_inst_req_1 : boolean;
  signal type_cast_376_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_390_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_390_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_390_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_390_inst_ack_1 : boolean;
  signal type_cast_394_inst_req_0 : boolean;
  signal type_cast_394_inst_ack_0 : boolean;
  signal type_cast_394_inst_req_1 : boolean;
  signal type_cast_394_inst_ack_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_408_inst_req_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_408_inst_ack_0 : boolean;
  signal RPIPE_Zeropad_input_pipe_408_inst_req_1 : boolean;
  signal RPIPE_Zeropad_input_pipe_408_inst_ack_1 : boolean;
  signal type_cast_412_inst_req_0 : boolean;
  signal type_cast_412_inst_ack_0 : boolean;
  signal type_cast_412_inst_req_1 : boolean;
  signal type_cast_412_inst_ack_1 : boolean;
  signal ptr_deref_420_store_0_req_0 : boolean;
  signal ptr_deref_420_store_0_ack_0 : boolean;
  signal ptr_deref_420_store_0_req_1 : boolean;
  signal ptr_deref_420_store_0_ack_1 : boolean;
  signal if_stmt_434_branch_req_0 : boolean;
  signal if_stmt_434_branch_ack_1 : boolean;
  signal if_stmt_434_branch_ack_0 : boolean;
  signal call_stmt_445_call_req_0 : boolean;
  signal call_stmt_445_call_ack_0 : boolean;
  signal call_stmt_445_call_req_1 : boolean;
  signal call_stmt_445_call_ack_1 : boolean;
  signal W_ifx_xthen191_exec_guard_823_delayed_1_0_856_inst_ack_0 : boolean;
  signal W_ifx_xthen191_exec_guard_823_delayed_1_0_856_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue208_exec_guard_863_delayed_1_0_917_inst_req_1 : boolean;
  signal phi_stmt_615_req_0 : boolean;
  signal W_landx_xlhsx_xtrue208_exec_guard_863_delayed_1_0_917_inst_ack_0 : boolean;
  signal W_landx_xlhsx_xtrue208_exec_guard_863_delayed_1_0_917_inst_req_0 : boolean;
  signal phi_stmt_615_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1451_inst_ack_0 : boolean;
  signal type_cast_854_inst_ack_1 : boolean;
  signal type_cast_854_inst_req_1 : boolean;
  signal phi_stmt_615_ack_0 : boolean;
  signal type_cast_854_inst_ack_0 : boolean;
  signal type_cast_854_inst_req_0 : boolean;
  signal type_cast_618_inst_req_0 : boolean;
  signal type_cast_618_inst_ack_0 : boolean;
  signal array_obj_ref_1187_index_offset_req_1 : boolean;
  signal type_cast_618_inst_req_1 : boolean;
  signal type_cast_618_inst_ack_1 : boolean;
  signal W_ifx_xthen180_exec_guard_768_delayed_6_0_792_inst_ack_1 : boolean;
  signal W_ifx_xthen180_exec_guard_768_delayed_6_0_792_inst_req_1 : boolean;
  signal W_output_byte_countx_x0_1017_delayed_2_0_1150_inst_ack_0 : boolean;
  signal type_cast_915_inst_ack_0 : boolean;
  signal MUX_842_inst_ack_1 : boolean;
  signal MUX_842_inst_req_1 : boolean;
  signal MUX_842_inst_ack_0 : boolean;
  signal MUX_842_inst_req_0 : boolean;
  signal type_cast_1210_inst_ack_0 : boolean;
  signal phi_stmt_620_req_0 : boolean;
  signal phi_stmt_620_req_1 : boolean;
  signal W_ifx_xthen180_ifx_xthen191_taken_807_delayed_12_0_833_inst_ack_1 : boolean;
  signal W_ifx_xthen180_ifx_xthen191_taken_807_delayed_12_0_833_inst_req_1 : boolean;
  signal phi_stmt_620_ack_0 : boolean;
  signal W_ifx_xthen180_ifx_xthen191_taken_807_delayed_12_0_833_inst_ack_0 : boolean;
  signal W_ifx_xthen180_ifx_xthen191_taken_807_delayed_12_0_833_inst_req_0 : boolean;
  signal type_cast_623_inst_req_0 : boolean;
  signal type_cast_623_inst_ack_0 : boolean;
  signal addr_of_790_final_reg_ack_0 : boolean;
  signal type_cast_623_inst_req_1 : boolean;
  signal type_cast_623_inst_ack_1 : boolean;
  signal MUX_1131_inst_req_1 : boolean;
  signal MUX_1131_inst_ack_1 : boolean;
  signal W_o1x_x1_860_delayed_1_0_909_inst_req_1 : boolean;
  signal type_cast_1210_inst_req_1 : boolean;
  signal W_o1x_x1_860_delayed_1_0_909_inst_ack_1 : boolean;
  signal phi_stmt_625_req_0 : boolean;
  signal W_output_byte_countx_x0_1017_delayed_2_0_1150_inst_req_1 : boolean;
  signal phi_stmt_625_req_1 : boolean;
  signal phi_stmt_625_ack_0 : boolean;
  signal addr_of_1188_final_reg_req_0 : boolean;
  signal addr_of_1188_final_reg_ack_0 : boolean;
  signal type_cast_628_inst_req_0 : boolean;
  signal type_cast_628_inst_ack_0 : boolean;
  signal type_cast_628_inst_req_1 : boolean;
  signal type_cast_628_inst_ack_1 : boolean;
  signal MUX_1099_inst_req_0 : boolean;
  signal W_output_byte_countx_x0_1017_delayed_2_0_1150_inst_ack_1 : boolean;
  signal type_cast_1470_inst_ack_0 : boolean;
  signal type_cast_1580_inst_ack_1 : boolean;
  signal addr_of_1188_final_reg_req_1 : boolean;
  signal phi_stmt_630_req_0 : boolean;
  signal addr_of_1188_final_reg_ack_1 : boolean;
  signal phi_stmt_630_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1436_inst_ack_1 : boolean;
  signal type_cast_1470_inst_ack_1 : boolean;
  signal phi_stmt_630_ack_0 : boolean;
  signal type_cast_633_inst_req_0 : boolean;
  signal type_cast_633_inst_ack_0 : boolean;
  signal type_cast_633_inst_req_1 : boolean;
  signal array_obj_ref_1521_index_offset_ack_0 : boolean;
  signal type_cast_633_inst_ack_1 : boolean;
  signal MUX_1099_inst_ack_0 : boolean;
  signal W_iNsTr_28_1010_delayed_2_0_1140_inst_req_0 : boolean;
  signal W_iNsTr_28_1010_delayed_2_0_1140_inst_ack_0 : boolean;
  signal type_cast_1470_inst_req_0 : boolean;
  signal phi_stmt_635_req_0 : boolean;
  signal MUX_1099_inst_req_1 : boolean;
  signal MUX_1099_inst_ack_1 : boolean;
  signal phi_stmt_635_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1436_inst_req_1 : boolean;
  signal phi_stmt_635_ack_0 : boolean;
  signal type_cast_1580_inst_req_1 : boolean;
  signal type_cast_638_inst_req_0 : boolean;
  signal type_cast_638_inst_ack_0 : boolean;
  signal type_cast_1530_inst_ack_0 : boolean;
  signal type_cast_638_inst_req_1 : boolean;
  signal type_cast_638_inst_ack_1 : boolean;
  signal ptr_deref_1192_store_0_req_1 : boolean;
  signal W_iNsTr_28_1010_delayed_2_0_1140_inst_req_1 : boolean;
  signal array_obj_ref_1521_index_offset_req_0 : boolean;
  signal W_iNsTr_28_1010_delayed_2_0_1140_inst_ack_1 : boolean;
  signal phi_stmt_640_req_0 : boolean;
  signal type_cast_1540_inst_ack_1 : boolean;
  signal phi_stmt_640_req_1 : boolean;
  signal phi_stmt_640_ack_0 : boolean;
  signal type_cast_643_inst_req_0 : boolean;
  signal type_cast_643_inst_ack_0 : boolean;
  signal type_cast_643_inst_req_1 : boolean;
  signal type_cast_643_inst_ack_1 : boolean;
  signal input_wordx_x1_at_entry_583_644_buf_req_0 : boolean;
  signal input_wordx_x1_at_entry_583_644_buf_ack_0 : boolean;
  signal input_wordx_x1_at_entry_583_644_buf_req_1 : boolean;
  signal input_wordx_x1_at_entry_583_644_buf_ack_1 : boolean;
  signal type_cast_684_inst_req_0 : boolean;
  signal type_cast_684_inst_ack_0 : boolean;
  signal type_cast_684_inst_req_1 : boolean;
  signal type_cast_684_inst_ack_1 : boolean;
  signal W_ifx_xend_exec_guard_686_delayed_1_0_686_inst_req_0 : boolean;
  signal W_ifx_xend_exec_guard_686_delayed_1_0_686_inst_ack_0 : boolean;
  signal W_ifx_xend_exec_guard_686_delayed_1_0_686_inst_req_1 : boolean;
  signal W_ifx_xend_exec_guard_686_delayed_1_0_686_inst_ack_1 : boolean;
  signal W_ifx_xend_exec_guard_693_delayed_1_0_696_inst_req_0 : boolean;
  signal W_ifx_xend_exec_guard_693_delayed_1_0_696_inst_ack_0 : boolean;
  signal W_ifx_xend_exec_guard_693_delayed_1_0_696_inst_req_1 : boolean;
  signal W_ifx_xend_exec_guard_693_delayed_1_0_696_inst_ack_1 : boolean;
  signal W_ifx_xend_exec_guard_700_delayed_1_0_706_inst_req_0 : boolean;
  signal W_ifx_xend_exec_guard_700_delayed_1_0_706_inst_ack_0 : boolean;
  signal W_ifx_xend_exec_guard_700_delayed_1_0_706_inst_req_1 : boolean;
  signal W_ifx_xend_exec_guard_700_delayed_1_0_706_inst_ack_1 : boolean;
  signal type_cast_712_inst_req_0 : boolean;
  signal type_cast_712_inst_ack_0 : boolean;
  signal type_cast_712_inst_req_1 : boolean;
  signal type_cast_712_inst_ack_1 : boolean;
  signal W_ifx_xend_exec_guard_705_delayed_2_0_714_inst_req_0 : boolean;
  signal W_ifx_xend_exec_guard_705_delayed_2_0_714_inst_ack_0 : boolean;
  signal W_ifx_xend_exec_guard_705_delayed_2_0_714_inst_req_1 : boolean;
  signal W_ifx_xend_exec_guard_705_delayed_2_0_714_inst_ack_1 : boolean;
  signal W_input_wordx_x1_707_delayed_2_0_717_inst_req_0 : boolean;
  signal W_input_wordx_x1_707_delayed_2_0_717_inst_ack_0 : boolean;
  signal W_input_wordx_x1_707_delayed_2_0_717_inst_req_1 : boolean;
  signal W_input_wordx_x1_707_delayed_2_0_717_inst_ack_1 : boolean;
  signal W_ifx_xend_exec_guard_718_delayed_2_0_733_inst_req_0 : boolean;
  signal W_ifx_xend_exec_guard_718_delayed_2_0_733_inst_ack_0 : boolean;
  signal W_ifx_xend_exec_guard_718_delayed_2_0_733_inst_req_1 : boolean;
  signal W_ifx_xend_exec_guard_718_delayed_2_0_733_inst_ack_1 : boolean;
  signal W_ifx_xend_exec_guard_725_delayed_2_0_743_inst_req_0 : boolean;
  signal W_ifx_xend_exec_guard_725_delayed_2_0_743_inst_ack_0 : boolean;
  signal W_ifx_xend_exec_guard_725_delayed_2_0_743_inst_req_1 : boolean;
  signal W_ifx_xend_exec_guard_725_delayed_2_0_743_inst_ack_1 : boolean;
  signal W_shl169_728_delayed_2_0_746_inst_req_0 : boolean;
  signal W_shl169_728_delayed_2_0_746_inst_ack_0 : boolean;
  signal W_shl169_728_delayed_2_0_746_inst_req_1 : boolean;
  signal W_shl169_728_delayed_2_0_746_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_926_inst_req_0 : boolean;
  signal type_cast_1210_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_926_inst_ack_0 : boolean;
  signal W_landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_926_inst_req_1 : boolean;
  signal W_landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_926_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1605_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1430_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1445_inst_ack_0 : boolean;
  signal array_obj_ref_1187_index_offset_ack_0 : boolean;
  signal array_obj_ref_1187_index_offset_req_0 : boolean;
  signal type_cast_1590_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_934_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_934_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1451_inst_req_1 : boolean;
  signal W_landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_934_inst_req_1 : boolean;
  signal W_landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_934_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1608_inst_req_0 : boolean;
  signal type_cast_1550_inst_req_0 : boolean;
  signal type_cast_1590_inst_ack_0 : boolean;
  signal W_o2x_x1_885_delayed_2_0_946_inst_req_0 : boolean;
  signal W_o2x_x1_885_delayed_2_0_946_inst_ack_0 : boolean;
  signal W_o2x_x1_885_delayed_2_0_946_inst_req_1 : boolean;
  signal W_o2x_x1_885_delayed_2_0_946_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1442_inst_req_0 : boolean;
  signal W_condx_xend_ifx_xend238_taken_997_delayed_1_0_1122_inst_ack_1 : boolean;
  signal type_cast_1590_inst_ack_1 : boolean;
  signal W_condx_xend_ifx_xend238_taken_997_delayed_1_0_1122_inst_req_1 : boolean;
  signal W_add_outx_x1_1059_delayed_2_0_1195_inst_ack_1 : boolean;
  signal W_add_outx_x1_1059_delayed_2_0_1195_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1451_inst_ack_1 : boolean;
  signal type_cast_952_inst_req_0 : boolean;
  signal type_cast_952_inst_ack_0 : boolean;
  signal type_cast_1091_inst_ack_0 : boolean;
  signal type_cast_952_inst_req_1 : boolean;
  signal type_cast_952_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1445_inst_req_1 : boolean;
  signal W_condx_xend_ifx_xend238_taken_997_delayed_1_0_1122_inst_ack_0 : boolean;
  signal type_cast_1091_inst_req_0 : boolean;
  signal W_target_out_offsetx_x1_890_delayed_2_0_954_inst_req_0 : boolean;
  signal W_add_outx_x1_1059_delayed_2_0_1195_inst_ack_0 : boolean;
  signal W_target_out_offsetx_x1_890_delayed_2_0_954_inst_ack_0 : boolean;
  signal W_target_out_offsetx_x1_890_delayed_2_0_954_inst_req_1 : boolean;
  signal W_add_outx_x1_1059_delayed_2_0_1195_inst_req_0 : boolean;
  signal W_target_out_offsetx_x1_890_delayed_2_0_954_inst_ack_1 : boolean;
  signal W_condx_xend_ifx_xend238_taken_997_delayed_1_0_1122_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1611_inst_ack_1 : boolean;
  signal type_cast_1540_inst_req_1 : boolean;
  signal W_landx_xlhsx_xtrue219_exec_guard_894_delayed_1_0_963_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue219_exec_guard_894_delayed_1_0_963_inst_ack_0 : boolean;
  signal W_landx_xlhsx_xtrue219_exec_guard_894_delayed_1_0_963_inst_req_1 : boolean;
  signal W_landx_xlhsx_xtrue219_exec_guard_894_delayed_1_0_963_inst_ack_1 : boolean;
  signal ptr_deref_1526_load_0_req_1 : boolean;
  signal type_cast_1470_inst_req_1 : boolean;
  signal W_landx_xlhsx_xtrue219_exec_guard_900_delayed_1_0_972_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue219_exec_guard_900_delayed_1_0_972_inst_ack_0 : boolean;
  signal W_landx_xlhsx_xtrue219_exec_guard_900_delayed_1_0_972_inst_req_1 : boolean;
  signal W_landx_xlhsx_xtrue219_exec_guard_900_delayed_1_0_972_inst_ack_1 : boolean;
  signal MUX_1113_inst_ack_1 : boolean;
  signal W_add234_903_delayed_1_0_975_inst_req_0 : boolean;
  signal W_add234_903_delayed_1_0_975_inst_ack_0 : boolean;
  signal type_cast_1590_inst_req_1 : boolean;
  signal W_add234_903_delayed_1_0_975_inst_req_1 : boolean;
  signal ptr_deref_1192_store_0_ack_1 : boolean;
  signal W_add234_903_delayed_1_0_975_inst_ack_1 : boolean;
  signal MUX_1113_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1445_inst_ack_1 : boolean;
  signal ptr_deref_1526_load_0_ack_1 : boolean;
  signal W_target_out_offsetx_x1_904_delayed_3_0_978_inst_req_0 : boolean;
  signal array_obj_ref_1521_index_offset_req_1 : boolean;
  signal W_target_out_offsetx_x1_904_delayed_3_0_978_inst_ack_0 : boolean;
  signal W_target_out_offsetx_x1_904_delayed_3_0_978_inst_req_1 : boolean;
  signal array_obj_ref_1521_index_offset_ack_1 : boolean;
  signal W_target_out_offsetx_x1_904_delayed_3_0_978_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1442_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1433_inst_req_0 : boolean;
  signal type_cast_1550_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1614_inst_ack_1 : boolean;
  signal W_ifx_xthen191_condx_xend_taken_911_delayed_1_0_991_inst_req_0 : boolean;
  signal W_ifx_xthen191_condx_xend_taken_911_delayed_1_0_991_inst_ack_0 : boolean;
  signal W_ifx_xthen191_condx_xend_taken_911_delayed_1_0_991_inst_req_1 : boolean;
  signal W_ifx_xthen191_condx_xend_taken_911_delayed_1_0_991_inst_ack_1 : boolean;
  signal W_ifx_xthen191_condx_xend_taken_918_delayed_2_0_1001_inst_req_0 : boolean;
  signal if_stmt_1461_branch_req_0 : boolean;
  signal W_ifx_xthen191_condx_xend_taken_918_delayed_2_0_1001_inst_ack_0 : boolean;
  signal W_ifx_xthen191_condx_xend_taken_918_delayed_2_0_1001_inst_req_1 : boolean;
  signal W_ifx_xthen191_condx_xend_taken_918_delayed_2_0_1001_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1442_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1442_inst_ack_1 : boolean;
  signal type_cast_1550_inst_req_1 : boolean;
  signal type_cast_1006_inst_req_0 : boolean;
  signal type_cast_1006_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1605_inst_req_1 : boolean;
  signal type_cast_1006_inst_req_1 : boolean;
  signal type_cast_1006_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1605_inst_ack_1 : boolean;
  signal type_cast_1550_inst_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue208_condx_xend_taken_921_delayed_1_0_1008_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue208_condx_xend_taken_921_delayed_1_0_1008_inst_ack_0 : boolean;
  signal W_landx_xlhsx_xtrue208_condx_xend_taken_921_delayed_1_0_1008_inst_req_1 : boolean;
  signal addr_of_1522_final_reg_req_0 : boolean;
  signal W_landx_xlhsx_xtrue208_condx_xend_taken_921_delayed_1_0_1008_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1433_inst_ack_0 : boolean;
  signal addr_of_1522_final_reg_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1433_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1433_inst_ack_1 : boolean;
  signal type_cast_1600_inst_req_0 : boolean;
  signal type_cast_1013_inst_req_0 : boolean;
  signal type_cast_1013_inst_ack_0 : boolean;
  signal type_cast_1013_inst_req_1 : boolean;
  signal type_cast_1013_inst_ack_1 : boolean;
  signal addr_of_1522_final_reg_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1439_inst_req_0 : boolean;
  signal W_landx_xlhsx_xtrue219_condx_xend_taken_924_delayed_1_0_1015_inst_req_0 : boolean;
  signal addr_of_1522_final_reg_ack_1 : boolean;
  signal W_landx_xlhsx_xtrue219_condx_xend_taken_924_delayed_1_0_1015_inst_ack_0 : boolean;
  signal type_cast_1600_inst_ack_0 : boolean;
  signal W_landx_xlhsx_xtrue219_condx_xend_taken_924_delayed_1_0_1015_inst_req_1 : boolean;
  signal W_landx_xlhsx_xtrue219_condx_xend_taken_924_delayed_1_0_1015_inst_ack_1 : boolean;
  signal if_stmt_1461_branch_ack_1 : boolean;
  signal W_condx_xend_exec_guard_933_delayed_1_0_1032_inst_req_0 : boolean;
  signal W_condx_xend_exec_guard_933_delayed_1_0_1032_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1439_inst_ack_0 : boolean;
  signal W_condx_xend_exec_guard_933_delayed_1_0_1032_inst_req_1 : boolean;
  signal W_condx_xend_exec_guard_933_delayed_1_0_1032_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1448_inst_req_0 : boolean;
  signal W_ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1045_inst_req_0 : boolean;
  signal W_ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1045_inst_ack_0 : boolean;
  signal W_ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1045_inst_req_1 : boolean;
  signal W_ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1045_inst_ack_1 : boolean;
  signal W_condx_xend_ifx_xend238_taken_949_delayed_10_0_1053_inst_req_0 : boolean;
  signal W_condx_xend_ifx_xend238_taken_949_delayed_10_0_1053_inst_ack_0 : boolean;
  signal W_condx_xend_ifx_xend238_taken_949_delayed_10_0_1053_inst_req_1 : boolean;
  signal W_condx_xend_ifx_xend238_taken_949_delayed_10_0_1053_inst_ack_1 : boolean;
  signal MUX_1062_inst_req_0 : boolean;
  signal MUX_1062_inst_ack_0 : boolean;
  signal MUX_1062_inst_req_1 : boolean;
  signal MUX_1062_inst_ack_1 : boolean;
  signal type_cast_1073_inst_req_0 : boolean;
  signal type_cast_1073_inst_ack_0 : boolean;
  signal type_cast_1073_inst_req_1 : boolean;
  signal type_cast_1073_inst_ack_1 : boolean;
  signal MUX_1081_inst_req_0 : boolean;
  signal MUX_1081_inst_ack_0 : boolean;
  signal MUX_1081_inst_req_1 : boolean;
  signal MUX_1081_inst_ack_1 : boolean;
  signal type_cast_1251_inst_req_0 : boolean;
  signal type_cast_1251_inst_ack_0 : boolean;
  signal type_cast_1251_inst_req_1 : boolean;
  signal type_cast_1251_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1614_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1614_inst_req_1 : boolean;
  signal ptr_deref_1526_load_0_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1451_inst_req_0 : boolean;
  signal ptr_deref_1526_load_0_req_0 : boolean;
  signal type_cast_1255_inst_req_0 : boolean;
  signal type_cast_1255_inst_ack_0 : boolean;
  signal type_cast_1580_inst_ack_0 : boolean;
  signal type_cast_1255_inst_req_1 : boolean;
  signal type_cast_1255_inst_ack_1 : boolean;
  signal type_cast_1580_inst_req_0 : boolean;
  signal type_cast_1271_inst_req_0 : boolean;
  signal type_cast_1271_inst_ack_0 : boolean;
  signal type_cast_1271_inst_req_1 : boolean;
  signal type_cast_1271_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1602_inst_ack_1 : boolean;
  signal W_o1x_x1_1134_delayed_2_0_1279_inst_req_0 : boolean;
  signal W_o1x_x1_1134_delayed_2_0_1279_inst_ack_0 : boolean;
  signal W_o1x_x1_1134_delayed_2_0_1279_inst_req_1 : boolean;
  signal W_o1x_x1_1134_delayed_2_0_1279_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1602_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1608_inst_ack_1 : boolean;
  signal W_inc265_1139_delayed_1_0_1287_inst_req_0 : boolean;
  signal W_inc265_1139_delayed_1_0_1287_inst_ack_0 : boolean;
  signal type_cast_1570_inst_ack_1 : boolean;
  signal W_inc265_1139_delayed_1_0_1287_inst_req_1 : boolean;
  signal W_inc265_1139_delayed_1_0_1287_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1602_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1611_inst_ack_0 : boolean;
  signal type_cast_1570_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1608_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1602_inst_req_0 : boolean;
  signal type_cast_1304_inst_req_0 : boolean;
  signal type_cast_1304_inst_ack_0 : boolean;
  signal type_cast_1570_inst_ack_0 : boolean;
  signal type_cast_1304_inst_req_1 : boolean;
  signal type_cast_1304_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1617_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1617_inst_ack_0 : boolean;
  signal type_cast_1540_inst_ack_0 : boolean;
  signal type_cast_1570_inst_req_0 : boolean;
  signal W_o0x_x1_1155_delayed_3_0_1306_inst_req_0 : boolean;
  signal W_o0x_x1_1155_delayed_3_0_1306_inst_ack_0 : boolean;
  signal W_o0x_x1_1155_delayed_3_0_1306_inst_req_1 : boolean;
  signal W_o0x_x1_1155_delayed_3_0_1306_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1614_inst_req_0 : boolean;
  signal type_cast_1540_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1611_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1617_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1617_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1608_inst_ack_0 : boolean;
  signal type_cast_1600_inst_ack_1 : boolean;
  signal do_while_stmt_588_branch_ack_0 : boolean;
  signal do_while_stmt_588_branch_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1436_inst_ack_0 : boolean;
  signal if_stmt_1332_branch_req_0 : boolean;
  signal type_cast_1600_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1436_inst_req_0 : boolean;
  signal if_stmt_1332_branch_ack_1 : boolean;
  signal if_stmt_1332_branch_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1611_inst_req_1 : boolean;
  signal type_cast_1560_inst_ack_1 : boolean;
  signal type_cast_1341_inst_req_0 : boolean;
  signal type_cast_1341_inst_ack_0 : boolean;
  signal type_cast_1560_inst_req_1 : boolean;
  signal type_cast_1341_inst_req_1 : boolean;
  signal type_cast_1479_inst_ack_1 : boolean;
  signal type_cast_1341_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1439_inst_ack_1 : boolean;
  signal type_cast_1479_inst_req_1 : boolean;
  signal call_stmt_1345_call_req_0 : boolean;
  signal call_stmt_1345_call_ack_0 : boolean;
  signal if_stmt_1461_branch_ack_0 : boolean;
  signal call_stmt_1345_call_req_1 : boolean;
  signal call_stmt_1345_call_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1439_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1448_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1448_inst_req_1 : boolean;
  signal type_cast_1530_inst_req_0 : boolean;
  signal type_cast_1479_inst_ack_0 : boolean;
  signal type_cast_1560_inst_ack_0 : boolean;
  signal type_cast_1349_inst_req_0 : boolean;
  signal type_cast_1479_inst_req_0 : boolean;
  signal type_cast_1349_inst_ack_0 : boolean;
  signal type_cast_1560_inst_req_0 : boolean;
  signal type_cast_1349_inst_req_1 : boolean;
  signal type_cast_1349_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1448_inst_ack_0 : boolean;
  signal type_cast_1358_inst_req_0 : boolean;
  signal type_cast_1358_inst_ack_0 : boolean;
  signal type_cast_1358_inst_req_1 : boolean;
  signal type_cast_1358_inst_ack_1 : boolean;
  signal type_cast_1368_inst_req_0 : boolean;
  signal type_cast_1368_inst_ack_0 : boolean;
  signal type_cast_1368_inst_req_1 : boolean;
  signal type_cast_1368_inst_ack_1 : boolean;
  signal type_cast_1378_inst_req_0 : boolean;
  signal type_cast_1378_inst_ack_0 : boolean;
  signal type_cast_1378_inst_req_1 : boolean;
  signal type_cast_1378_inst_ack_1 : boolean;
  signal type_cast_1388_inst_req_0 : boolean;
  signal type_cast_1388_inst_ack_0 : boolean;
  signal type_cast_1388_inst_req_1 : boolean;
  signal type_cast_1388_inst_ack_1 : boolean;
  signal type_cast_1398_inst_req_0 : boolean;
  signal type_cast_1398_inst_ack_0 : boolean;
  signal type_cast_1398_inst_req_1 : boolean;
  signal type_cast_1398_inst_ack_1 : boolean;
  signal type_cast_1408_inst_req_0 : boolean;
  signal type_cast_1408_inst_ack_0 : boolean;
  signal type_cast_1408_inst_req_1 : boolean;
  signal type_cast_1408_inst_ack_1 : boolean;
  signal type_cast_1418_inst_req_0 : boolean;
  signal type_cast_1418_inst_ack_0 : boolean;
  signal type_cast_1418_inst_req_1 : boolean;
  signal type_cast_1418_inst_ack_1 : boolean;
  signal type_cast_1428_inst_req_0 : boolean;
  signal type_cast_1428_inst_ack_0 : boolean;
  signal type_cast_1428_inst_req_1 : boolean;
  signal type_cast_1428_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1430_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1430_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1620_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1620_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1620_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1620_inst_ack_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1623_inst_req_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1623_inst_ack_0 : boolean;
  signal WPIPE_Zeropad_output_pipe_1623_inst_req_1 : boolean;
  signal WPIPE_Zeropad_output_pipe_1623_inst_ack_1 : boolean;
  signal if_stmt_1637_branch_req_0 : boolean;
  signal if_stmt_1637_branch_ack_1 : boolean;
  signal if_stmt_1637_branch_ack_0 : boolean;
  signal phi_stmt_269_req_0 : boolean;
  signal type_cast_275_inst_req_0 : boolean;
  signal type_cast_275_inst_ack_0 : boolean;
  signal type_cast_275_inst_req_1 : boolean;
  signal type_cast_275_inst_ack_1 : boolean;
  signal phi_stmt_269_req_1 : boolean;
  signal phi_stmt_269_ack_0 : boolean;
  signal type_cast_542_inst_req_0 : boolean;
  signal type_cast_542_inst_ack_0 : boolean;
  signal type_cast_542_inst_req_1 : boolean;
  signal type_cast_542_inst_ack_1 : boolean;
  signal phi_stmt_539_req_0 : boolean;
  signal type_cast_586_inst_req_0 : boolean;
  signal type_cast_586_inst_ack_0 : boolean;
  signal type_cast_586_inst_req_1 : boolean;
  signal type_cast_586_inst_ack_1 : boolean;
  signal phi_stmt_583_req_0 : boolean;
  signal phi_stmt_539_ack_0 : boolean;
  signal phi_stmt_583_ack_0 : boolean;
  signal phi_stmt_1507_req_0 : boolean;
  signal type_cast_1513_inst_req_0 : boolean;
  signal type_cast_1513_inst_ack_0 : boolean;
  signal type_cast_1513_inst_req_1 : boolean;
  signal type_cast_1513_inst_ack_1 : boolean;
  signal phi_stmt_1507_req_1 : boolean;
  signal phi_stmt_1507_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad_CP_182_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad_CP_182_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad_CP_182_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad_CP_182_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad_CP_182: Block -- control-path 
    signal zeropad_CP_182_elements: BooleanArray(740 downto 0);
    -- 
  begin -- 
    zeropad_CP_182_elements(0) <= zeropad_CP_182_start;
    zeropad_CP_182_symbol <= zeropad_CP_182_elements(740);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	25 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	29 
    -- CP-element group 0: 	33 
    -- CP-element group 0: 	37 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	45 
    -- CP-element group 0: 	49 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	55 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (50) 
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_63_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_43/$entry
      -- CP-element group 0: 	 branch_block_stmt_43/branch_block_stmt_43__entry__
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230__entry__
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/$entry
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_45_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_45_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_45_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_50_update_start_
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_50_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_50_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_63_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_63_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_75_update_start_
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_75_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_75_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_88_update_start_
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_88_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_88_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_100_update_start_
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_100_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_100_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_113_update_start_
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_113_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_113_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_126_update_start_
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_126_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_126_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_139_update_start_
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_139_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_139_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_151_update_start_
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_151_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_151_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_164_update_start_
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_164_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_164_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_176_update_start_
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_176_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_176_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_189_update_start_
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_189_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_189_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_208_update_start_
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_208_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_208_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_212_update_start_
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_212_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_212_Update/cr
      -- 
    rr_254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(0), ack => RPIPE_Zeropad_input_pipe_45_inst_req_0); -- 
    cr_273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(0), ack => type_cast_50_inst_req_1); -- 
    cr_301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(0), ack => type_cast_63_inst_req_1); -- 
    cr_329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(0), ack => type_cast_75_inst_req_1); -- 
    cr_357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(0), ack => type_cast_88_inst_req_1); -- 
    cr_385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(0), ack => type_cast_100_inst_req_1); -- 
    cr_413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(0), ack => type_cast_113_inst_req_1); -- 
    cr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(0), ack => type_cast_126_inst_req_1); -- 
    cr_469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(0), ack => type_cast_139_inst_req_1); -- 
    cr_497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(0), ack => type_cast_151_inst_req_1); -- 
    cr_525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(0), ack => type_cast_164_inst_req_1); -- 
    cr_553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(0), ack => type_cast_176_inst_req_1); -- 
    cr_581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(0), ack => type_cast_189_inst_req_1); -- 
    cr_595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(0), ack => type_cast_208_inst_req_1); -- 
    cr_609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(0), ack => type_cast_212_inst_req_1); -- 
    -- CP-element group 1:  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	614 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	615 
    -- CP-element group 1: 	616 
    -- CP-element group 1:  members (9) 
      -- CP-element group 1: 	 branch_block_stmt_43/do_while_stmt_588__exit__
      -- CP-element group 1: 	 branch_block_stmt_43/if_stmt_1332__entry__
      -- CP-element group 1: 	 branch_block_stmt_43/if_stmt_1332_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_43/if_stmt_1332_eval_test/$entry
      -- CP-element group 1: 	 branch_block_stmt_43/if_stmt_1332_eval_test/$exit
      -- CP-element group 1: 	 branch_block_stmt_43/if_stmt_1332_eval_test/branch_req
      -- CP-element group 1: 	 branch_block_stmt_43/R_ifx_xend253_whilex_xend_taken_1333_place
      -- CP-element group 1: 	 branch_block_stmt_43/if_stmt_1332_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_43/if_stmt_1332_else_link/$entry
      -- 
    branch_req_2620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(1), ack => if_stmt_1332_branch_req_0); -- 
    zeropad_CP_182_elements(1) <= zeropad_CP_182_elements(614);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_45_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_45_update_start_
      -- CP-element group 2: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_45_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_45_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_45_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_45_Update/cr
      -- 
    ra_255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_45_inst_ack_0, ack => zeropad_CP_182_elements(2)); -- 
    cr_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(2), ack => RPIPE_Zeropad_input_pipe_45_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	6 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_59_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_45_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_45_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_45_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_50_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_50_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_50_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_59_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_59_Sample/$entry
      -- 
    ca_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_45_inst_ack_1, ack => zeropad_CP_182_elements(3)); -- 
    rr_282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(3), ack => RPIPE_Zeropad_input_pipe_59_inst_req_0); -- 
    rr_268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(3), ack => type_cast_50_inst_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_50_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_50_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_50_Sample/ra
      -- 
    ra_269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_50_inst_ack_0, ack => zeropad_CP_182_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	56 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_50_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_50_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_50_Update/ca
      -- 
    ca_274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_50_inst_ack_1, ack => zeropad_CP_182_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_59_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_59_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_59_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_59_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_59_update_start_
      -- CP-element group 6: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_59_Sample/$exit
      -- 
    ra_283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_59_inst_ack_0, ack => zeropad_CP_182_elements(6)); -- 
    cr_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(6), ack => RPIPE_Zeropad_input_pipe_59_inst_req_1); -- 
    -- CP-element group 7:  fork  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	10 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_59_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_59_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_63_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_59_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_63_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_63_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_71_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_71_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_71_Sample/rr
      -- 
    ca_288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_59_inst_ack_1, ack => zeropad_CP_182_elements(7)); -- 
    rr_296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(7), ack => type_cast_63_inst_req_0); -- 
    rr_310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(7), ack => RPIPE_Zeropad_input_pipe_71_inst_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_63_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_63_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_63_Sample/ra
      -- 
    ra_297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_0, ack => zeropad_CP_182_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	56 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_63_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_63_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_63_Update/ca
      -- 
    ca_302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_1, ack => zeropad_CP_182_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	7 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_71_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_71_update_start_
      -- CP-element group 10: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_71_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_71_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_71_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_71_Update/cr
      -- 
    ra_311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_71_inst_ack_0, ack => zeropad_CP_182_elements(10)); -- 
    cr_315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(10), ack => RPIPE_Zeropad_input_pipe_71_inst_req_1); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_71_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_71_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_71_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_75_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_75_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_75_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_84_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_84_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_84_Sample/rr
      -- 
    ca_316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_71_inst_ack_1, ack => zeropad_CP_182_elements(11)); -- 
    rr_324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(11), ack => type_cast_75_inst_req_0); -- 
    rr_338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(11), ack => RPIPE_Zeropad_input_pipe_84_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_75_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_75_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_75_Sample/ra
      -- 
    ra_325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_75_inst_ack_0, ack => zeropad_CP_182_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	56 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_75_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_75_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_75_Update/ca
      -- 
    ca_330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_75_inst_ack_1, ack => zeropad_CP_182_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_84_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_84_update_start_
      -- CP-element group 14: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_84_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_84_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_84_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_84_Update/cr
      -- 
    ra_339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_84_inst_ack_0, ack => zeropad_CP_182_elements(14)); -- 
    cr_343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(14), ack => RPIPE_Zeropad_input_pipe_84_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	18 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_84_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_84_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_84_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_88_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_88_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_88_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_96_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_96_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_96_Sample/rr
      -- 
    ca_344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_84_inst_ack_1, ack => zeropad_CP_182_elements(15)); -- 
    rr_352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(15), ack => type_cast_88_inst_req_0); -- 
    rr_366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(15), ack => RPIPE_Zeropad_input_pipe_96_inst_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_88_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_88_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_88_Sample/ra
      -- 
    ra_353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_88_inst_ack_0, ack => zeropad_CP_182_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	56 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_88_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_88_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_88_Update/ca
      -- 
    ca_358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_88_inst_ack_1, ack => zeropad_CP_182_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_96_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_96_update_start_
      -- CP-element group 18: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_96_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_96_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_96_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_96_Update/cr
      -- 
    ra_367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_96_inst_ack_0, ack => zeropad_CP_182_elements(18)); -- 
    cr_371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(18), ack => RPIPE_Zeropad_input_pipe_96_inst_req_1); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_96_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_96_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_96_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_100_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_100_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_100_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_109_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_109_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_109_Sample/rr
      -- 
    ca_372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_96_inst_ack_1, ack => zeropad_CP_182_elements(19)); -- 
    rr_380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(19), ack => type_cast_100_inst_req_0); -- 
    rr_394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(19), ack => RPIPE_Zeropad_input_pipe_109_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_100_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_100_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_100_Sample/ra
      -- 
    ra_381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_100_inst_ack_0, ack => zeropad_CP_182_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	56 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_100_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_100_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_100_Update/ca
      -- 
    ca_386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_100_inst_ack_1, ack => zeropad_CP_182_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_109_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_109_update_start_
      -- CP-element group 22: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_109_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_109_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_109_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_109_Update/cr
      -- 
    ra_395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_109_inst_ack_0, ack => zeropad_CP_182_elements(22)); -- 
    cr_399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(22), ack => RPIPE_Zeropad_input_pipe_109_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	26 
    -- CP-element group 23:  members (9) 
      -- CP-element group 23: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_109_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_109_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_109_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_113_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_113_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_113_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_121_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_121_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_121_Sample/rr
      -- 
    ca_400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_109_inst_ack_1, ack => zeropad_CP_182_elements(23)); -- 
    rr_408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(23), ack => type_cast_113_inst_req_0); -- 
    rr_422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(23), ack => RPIPE_Zeropad_input_pipe_121_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_113_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_113_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_113_Sample/ra
      -- 
    ra_409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_113_inst_ack_0, ack => zeropad_CP_182_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	0 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	56 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_113_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_113_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_113_Update/ca
      -- 
    ca_414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_113_inst_ack_1, ack => zeropad_CP_182_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	23 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_121_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_121_update_start_
      -- CP-element group 26: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_121_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_121_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_121_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_121_Update/cr
      -- 
    ra_423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_121_inst_ack_0, ack => zeropad_CP_182_elements(26)); -- 
    cr_427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(26), ack => RPIPE_Zeropad_input_pipe_121_inst_req_1); -- 
    -- CP-element group 27:  fork  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	30 
    -- CP-element group 27:  members (9) 
      -- CP-element group 27: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_121_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_121_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_121_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_126_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_126_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_126_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_135_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_135_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_135_Sample/rr
      -- 
    ca_428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_121_inst_ack_1, ack => zeropad_CP_182_elements(27)); -- 
    rr_436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(27), ack => type_cast_126_inst_req_0); -- 
    rr_450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(27), ack => RPIPE_Zeropad_input_pipe_135_inst_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_126_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_126_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_126_Sample/ra
      -- 
    ra_437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_0, ack => zeropad_CP_182_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	0 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	50 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_126_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_126_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_126_Update/ca
      -- 
    ca_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_1, ack => zeropad_CP_182_elements(29)); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_135_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_135_update_start_
      -- CP-element group 30: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_135_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_135_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_135_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_135_Update/cr
      -- 
    ra_451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_135_inst_ack_0, ack => zeropad_CP_182_elements(30)); -- 
    cr_455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(30), ack => RPIPE_Zeropad_input_pipe_135_inst_req_1); -- 
    -- CP-element group 31:  fork  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_135_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_135_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_135_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_139_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_139_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_139_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_147_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_147_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_147_Sample/rr
      -- 
    ca_456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_135_inst_ack_1, ack => zeropad_CP_182_elements(31)); -- 
    rr_464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(31), ack => type_cast_139_inst_req_0); -- 
    rr_478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(31), ack => RPIPE_Zeropad_input_pipe_147_inst_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_139_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_139_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_139_Sample/ra
      -- 
    ra_465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_139_inst_ack_0, ack => zeropad_CP_182_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	50 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_139_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_139_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_139_Update/ca
      -- 
    ca_470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_139_inst_ack_1, ack => zeropad_CP_182_elements(33)); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_147_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_147_update_start_
      -- CP-element group 34: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_147_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_147_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_147_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_147_Update/cr
      -- 
    ra_479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_147_inst_ack_0, ack => zeropad_CP_182_elements(34)); -- 
    cr_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(34), ack => RPIPE_Zeropad_input_pipe_147_inst_req_1); -- 
    -- CP-element group 35:  fork  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (9) 
      -- CP-element group 35: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_147_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_147_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_147_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_151_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_151_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_151_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_160_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_160_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_160_Sample/rr
      -- 
    ca_484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_147_inst_ack_1, ack => zeropad_CP_182_elements(35)); -- 
    rr_492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(35), ack => type_cast_151_inst_req_0); -- 
    rr_506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(35), ack => RPIPE_Zeropad_input_pipe_160_inst_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_151_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_151_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_151_Sample/ra
      -- 
    ra_493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_151_inst_ack_0, ack => zeropad_CP_182_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	0 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	53 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_151_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_151_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_151_Update/ca
      -- 
    ca_498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_151_inst_ack_1, ack => zeropad_CP_182_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_160_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_160_update_start_
      -- CP-element group 38: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_160_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_160_Sample/ra
      -- CP-element group 38: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_160_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_160_Update/cr
      -- 
    ra_507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_160_inst_ack_0, ack => zeropad_CP_182_elements(38)); -- 
    cr_511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(38), ack => RPIPE_Zeropad_input_pipe_160_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39: 	42 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_160_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_160_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_160_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_164_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_164_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_164_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_172_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_172_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_172_Sample/rr
      -- 
    ca_512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_160_inst_ack_1, ack => zeropad_CP_182_elements(39)); -- 
    rr_520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(39), ack => type_cast_164_inst_req_0); -- 
    rr_534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(39), ack => RPIPE_Zeropad_input_pipe_172_inst_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_164_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_164_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_164_Sample/ra
      -- 
    ra_521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_164_inst_ack_0, ack => zeropad_CP_182_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	53 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_164_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_164_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_164_Update/ca
      -- 
    ca_526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_164_inst_ack_1, ack => zeropad_CP_182_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	39 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_172_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_172_update_start_
      -- CP-element group 42: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_172_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_172_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_172_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_172_Update/cr
      -- 
    ra_535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_172_inst_ack_0, ack => zeropad_CP_182_elements(42)); -- 
    cr_539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(42), ack => RPIPE_Zeropad_input_pipe_172_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43: 	46 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_172_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_172_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_172_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_176_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_176_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_176_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_185_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_185_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_185_Sample/rr
      -- 
    ca_540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_172_inst_ack_1, ack => zeropad_CP_182_elements(43)); -- 
    rr_548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(43), ack => type_cast_176_inst_req_0); -- 
    rr_562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(43), ack => RPIPE_Zeropad_input_pipe_185_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_176_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_176_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_176_Sample/ra
      -- 
    ra_549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_176_inst_ack_0, ack => zeropad_CP_182_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	0 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	56 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_176_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_176_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_176_Update/ca
      -- 
    ca_554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_176_inst_ack_1, ack => zeropad_CP_182_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	43 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_185_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_185_update_start_
      -- CP-element group 46: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_185_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_185_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_185_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_185_Update/cr
      -- 
    ra_563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_185_inst_ack_0, ack => zeropad_CP_182_elements(46)); -- 
    cr_567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(46), ack => RPIPE_Zeropad_input_pipe_185_inst_req_1); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_185_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_185_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/RPIPE_Zeropad_input_pipe_185_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_189_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_189_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_189_Sample/rr
      -- 
    ca_568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_185_inst_ack_1, ack => zeropad_CP_182_elements(47)); -- 
    rr_576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(47), ack => type_cast_189_inst_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_189_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_189_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_189_Sample/ra
      -- 
    ra_577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_189_inst_ack_0, ack => zeropad_CP_182_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	0 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	56 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_189_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_189_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_189_Update/ca
      -- 
    ca_582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_189_inst_ack_1, ack => zeropad_CP_182_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	29 
    -- CP-element group 50: 	33 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_208_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_208_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_208_Sample/rr
      -- 
    rr_590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(50), ack => type_cast_208_inst_req_0); -- 
    zeropad_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "zeropad_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(29) & zeropad_CP_182_elements(33);
      gj_zeropad_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_208_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_208_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_208_Sample/ra
      -- 
    ra_591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_208_inst_ack_0, ack => zeropad_CP_182_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	56 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_208_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_208_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_208_Update/ca
      -- 
    ca_596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_208_inst_ack_1, ack => zeropad_CP_182_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	37 
    -- CP-element group 53: 	41 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_212_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_212_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_212_Sample/rr
      -- 
    rr_604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(53), ack => type_cast_212_inst_req_0); -- 
    zeropad_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "zeropad_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(37) & zeropad_CP_182_elements(41);
      gj_zeropad_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_212_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_212_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_212_Sample/ra
      -- 
    ra_605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_212_inst_ack_0, ack => zeropad_CP_182_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	0 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_212_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_212_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/type_cast_212_Update/ca
      -- 
    ca_610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_212_inst_ack_1, ack => zeropad_CP_182_elements(55)); -- 
    -- CP-element group 56:  branch  join  transition  place  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	9 
    -- CP-element group 56: 	13 
    -- CP-element group 56: 	17 
    -- CP-element group 56: 	21 
    -- CP-element group 56: 	25 
    -- CP-element group 56: 	5 
    -- CP-element group 56: 	45 
    -- CP-element group 56: 	49 
    -- CP-element group 56: 	52 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (10) 
      -- CP-element group 56: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230__exit__
      -- CP-element group 56: 	 branch_block_stmt_43/if_stmt_231__entry__
      -- CP-element group 56: 	 branch_block_stmt_43/assign_stmt_46_to_assign_stmt_230/$exit
      -- CP-element group 56: 	 branch_block_stmt_43/if_stmt_231_dead_link/$entry
      -- CP-element group 56: 	 branch_block_stmt_43/if_stmt_231_eval_test/$entry
      -- CP-element group 56: 	 branch_block_stmt_43/if_stmt_231_eval_test/$exit
      -- CP-element group 56: 	 branch_block_stmt_43/if_stmt_231_eval_test/branch_req
      -- CP-element group 56: 	 branch_block_stmt_43/R_cmp462_232_place
      -- CP-element group 56: 	 branch_block_stmt_43/if_stmt_231_if_link/$entry
      -- CP-element group 56: 	 branch_block_stmt_43/if_stmt_231_else_link/$entry
      -- 
    branch_req_618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(56), ack => if_stmt_231_branch_req_0); -- 
    zeropad_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 27) := "zeropad_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(9) & zeropad_CP_182_elements(13) & zeropad_CP_182_elements(17) & zeropad_CP_182_elements(21) & zeropad_CP_182_elements(25) & zeropad_CP_182_elements(5) & zeropad_CP_182_elements(45) & zeropad_CP_182_elements(49) & zeropad_CP_182_elements(52) & zeropad_CP_182_elements(55);
      gj_zeropad_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  merge  transition  place  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	717 
    -- CP-element group 57:  members (18) 
      -- CP-element group 57: 	 branch_block_stmt_43/merge_stmt_237__exit__
      -- CP-element group 57: 	 branch_block_stmt_43/assign_stmt_242_to_assign_stmt_266__entry__
      -- CP-element group 57: 	 branch_block_stmt_43/assign_stmt_242_to_assign_stmt_266__exit__
      -- CP-element group 57: 	 branch_block_stmt_43/bbx_xnph464_forx_xbody
      -- CP-element group 57: 	 branch_block_stmt_43/if_stmt_231_if_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_43/if_stmt_231_if_link/if_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_43/entry_bbx_xnph464
      -- CP-element group 57: 	 branch_block_stmt_43/assign_stmt_242_to_assign_stmt_266/$entry
      -- CP-element group 57: 	 branch_block_stmt_43/assign_stmt_242_to_assign_stmt_266/$exit
      -- CP-element group 57: 	 branch_block_stmt_43/entry_bbx_xnph464_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_43/entry_bbx_xnph464_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_43/merge_stmt_237_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_43/merge_stmt_237_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_43/merge_stmt_237_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_43/merge_stmt_237_PhiAck/dummy
      -- CP-element group 57: 	 branch_block_stmt_43/bbx_xnph464_forx_xbody_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_43/bbx_xnph464_forx_xbody_PhiReq/phi_stmt_269/$entry
      -- CP-element group 57: 	 branch_block_stmt_43/bbx_xnph464_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_sources/$entry
      -- 
    if_choice_transition_623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_231_branch_ack_1, ack => zeropad_CP_182_elements(57)); -- 
    -- CP-element group 58:  transition  place  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	723 
    -- CP-element group 58:  members (5) 
      -- CP-element group 58: 	 branch_block_stmt_43/if_stmt_231_else_link/$exit
      -- CP-element group 58: 	 branch_block_stmt_43/if_stmt_231_else_link/else_choice_transition
      -- CP-element group 58: 	 branch_block_stmt_43/entry_forx_xend
      -- CP-element group 58: 	 branch_block_stmt_43/entry_forx_xend_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_43/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_231_branch_ack_0, ack => zeropad_CP_182_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	722 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	98 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_final_index_sum_regn_sample_complete
      -- CP-element group 59: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_final_index_sum_regn_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_final_index_sum_regn_Sample/ack
      -- 
    ack_661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_283_index_offset_ack_0, ack => zeropad_CP_182_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	722 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (11) 
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/addr_of_284_request/$entry
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/addr_of_284_request/req
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/addr_of_284_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_root_address_calculated
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_offset_calculated
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_final_index_sum_regn_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_final_index_sum_regn_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_base_plus_offset/$entry
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_base_plus_offset/$exit
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_base_plus_offset/sum_rename_req
      -- CP-element group 60: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_base_plus_offset/sum_rename_ack
      -- 
    ack_666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_283_index_offset_ack_1, ack => zeropad_CP_182_elements(60)); -- 
    req_675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(60), ack => addr_of_284_final_reg_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/addr_of_284_request/$exit
      -- CP-element group 61: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/addr_of_284_request/ack
      -- CP-element group 61: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/addr_of_284_sample_completed_
      -- 
    ack_676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_284_final_reg_ack_0, ack => zeropad_CP_182_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	722 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	95 
    -- CP-element group 62:  members (19) 
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/addr_of_284_complete/$exit
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/addr_of_284_complete/ack
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/addr_of_284_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_base_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_word_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_root_address_calculated
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_base_address_resized
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_base_addr_resize/$entry
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_base_addr_resize/$exit
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_base_addr_resize/base_resize_req
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_base_addr_resize/base_resize_ack
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_base_plus_offset/$entry
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_base_plus_offset/$exit
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_base_plus_offset/sum_rename_req
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_base_plus_offset/sum_rename_ack
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_word_addrgen/$entry
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_word_addrgen/$exit
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_word_addrgen/root_register_req
      -- CP-element group 62: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_word_addrgen/root_register_ack
      -- 
    ack_681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_284_final_reg_ack_1, ack => zeropad_CP_182_elements(62)); -- 
    -- CP-element group 63:  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	722 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_287_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_287_update_start_
      -- CP-element group 63: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_287_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_287_Sample/ra
      -- CP-element group 63: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_287_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_287_Update/cr
      -- 
    ra_690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_287_inst_ack_0, ack => zeropad_CP_182_elements(63)); -- 
    cr_694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(63), ack => RPIPE_Zeropad_input_pipe_287_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: 	67 
    -- CP-element group 64:  members (9) 
      -- CP-element group 64: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_287_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_287_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_287_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_291_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_291_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_291_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_300_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_300_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_300_Sample/rr
      -- 
    ca_695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_287_inst_ack_1, ack => zeropad_CP_182_elements(64)); -- 
    rr_703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(64), ack => type_cast_291_inst_req_0); -- 
    rr_717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(64), ack => RPIPE_Zeropad_input_pipe_300_inst_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_291_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_291_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_291_Sample/ra
      -- 
    ra_704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_291_inst_ack_0, ack => zeropad_CP_182_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	722 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	95 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_291_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_291_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_291_Update/ca
      -- 
    ca_709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_291_inst_ack_1, ack => zeropad_CP_182_elements(66)); -- 
    -- CP-element group 67:  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	64 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (6) 
      -- CP-element group 67: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_300_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_300_update_start_
      -- CP-element group 67: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_300_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_300_Sample/ra
      -- CP-element group 67: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_300_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_300_Update/cr
      -- 
    ra_718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_300_inst_ack_0, ack => zeropad_CP_182_elements(67)); -- 
    cr_722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(67), ack => RPIPE_Zeropad_input_pipe_300_inst_req_1); -- 
    -- CP-element group 68:  fork  transition  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	71 
    -- CP-element group 68:  members (9) 
      -- CP-element group 68: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_300_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_300_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_300_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_304_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_304_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_304_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_318_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_318_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_318_Sample/rr
      -- 
    ca_723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_300_inst_ack_1, ack => zeropad_CP_182_elements(68)); -- 
    rr_731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(68), ack => type_cast_304_inst_req_0); -- 
    rr_745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(68), ack => RPIPE_Zeropad_input_pipe_318_inst_req_0); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_304_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_304_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_304_Sample/ra
      -- 
    ra_732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_304_inst_ack_0, ack => zeropad_CP_182_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	722 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	95 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_304_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_304_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_304_Update/ca
      -- 
    ca_737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_304_inst_ack_1, ack => zeropad_CP_182_elements(70)); -- 
    -- CP-element group 71:  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	68 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (6) 
      -- CP-element group 71: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_318_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_318_update_start_
      -- CP-element group 71: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_318_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_318_Sample/ra
      -- CP-element group 71: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_318_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_318_Update/cr
      -- 
    ra_746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_318_inst_ack_0, ack => zeropad_CP_182_elements(71)); -- 
    cr_750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(71), ack => RPIPE_Zeropad_input_pipe_318_inst_req_1); -- 
    -- CP-element group 72:  fork  transition  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72: 	75 
    -- CP-element group 72:  members (9) 
      -- CP-element group 72: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_318_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_318_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_318_Update/ca
      -- CP-element group 72: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_322_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_322_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_322_Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_336_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_336_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_336_Sample/rr
      -- 
    ca_751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_318_inst_ack_1, ack => zeropad_CP_182_elements(72)); -- 
    rr_759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(72), ack => type_cast_322_inst_req_0); -- 
    rr_773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(72), ack => RPIPE_Zeropad_input_pipe_336_inst_req_0); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_322_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_322_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_322_Sample/ra
      -- 
    ra_760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_322_inst_ack_0, ack => zeropad_CP_182_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	722 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	95 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_322_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_322_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_322_Update/ca
      -- 
    ca_765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_322_inst_ack_1, ack => zeropad_CP_182_elements(74)); -- 
    -- CP-element group 75:  transition  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	72 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (6) 
      -- CP-element group 75: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_336_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_336_update_start_
      -- CP-element group 75: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_336_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_336_Sample/ra
      -- CP-element group 75: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_336_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_336_Update/cr
      -- 
    ra_774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_336_inst_ack_0, ack => zeropad_CP_182_elements(75)); -- 
    cr_778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(75), ack => RPIPE_Zeropad_input_pipe_336_inst_req_1); -- 
    -- CP-element group 76:  fork  transition  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	79 
    -- CP-element group 76:  members (9) 
      -- CP-element group 76: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_336_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_336_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_336_Update/ca
      -- CP-element group 76: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_340_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_340_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_340_Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_354_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_354_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_354_Sample/rr
      -- 
    ca_779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_336_inst_ack_1, ack => zeropad_CP_182_elements(76)); -- 
    rr_787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(76), ack => type_cast_340_inst_req_0); -- 
    rr_801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(76), ack => RPIPE_Zeropad_input_pipe_354_inst_req_0); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_340_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_340_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_340_Sample/ra
      -- 
    ra_788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_340_inst_ack_0, ack => zeropad_CP_182_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	722 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	95 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_340_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_340_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_340_Update/ca
      -- 
    ca_793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_340_inst_ack_1, ack => zeropad_CP_182_elements(78)); -- 
    -- CP-element group 79:  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	76 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (6) 
      -- CP-element group 79: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_354_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_354_update_start_
      -- CP-element group 79: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_354_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_354_Sample/ra
      -- CP-element group 79: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_354_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_354_Update/cr
      -- 
    ra_802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_354_inst_ack_0, ack => zeropad_CP_182_elements(79)); -- 
    cr_806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(79), ack => RPIPE_Zeropad_input_pipe_354_inst_req_1); -- 
    -- CP-element group 80:  fork  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (9) 
      -- CP-element group 80: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_354_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_354_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_354_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_358_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_358_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_358_Sample/rr
      -- CP-element group 80: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_372_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_372_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_372_Sample/rr
      -- 
    ca_807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_354_inst_ack_1, ack => zeropad_CP_182_elements(80)); -- 
    rr_815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(80), ack => type_cast_358_inst_req_0); -- 
    rr_829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(80), ack => RPIPE_Zeropad_input_pipe_372_inst_req_0); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_358_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_358_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_358_Sample/ra
      -- 
    ra_816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_358_inst_ack_0, ack => zeropad_CP_182_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	722 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	95 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_358_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_358_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_358_Update/ca
      -- 
    ca_821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_358_inst_ack_1, ack => zeropad_CP_182_elements(82)); -- 
    -- CP-element group 83:  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	80 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (6) 
      -- CP-element group 83: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_372_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_372_update_start_
      -- CP-element group 83: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_372_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_372_Sample/ra
      -- CP-element group 83: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_372_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_372_Update/cr
      -- 
    ra_830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_372_inst_ack_0, ack => zeropad_CP_182_elements(83)); -- 
    cr_834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(83), ack => RPIPE_Zeropad_input_pipe_372_inst_req_1); -- 
    -- CP-element group 84:  fork  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84: 	87 
    -- CP-element group 84:  members (9) 
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_372_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_372_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_372_Update/ca
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_376_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_376_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_376_Sample/rr
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_390_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_390_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_390_Sample/rr
      -- 
    ca_835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_372_inst_ack_1, ack => zeropad_CP_182_elements(84)); -- 
    rr_843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(84), ack => type_cast_376_inst_req_0); -- 
    rr_857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(84), ack => RPIPE_Zeropad_input_pipe_390_inst_req_0); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_376_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_376_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_376_Sample/ra
      -- 
    ra_844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_376_inst_ack_0, ack => zeropad_CP_182_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	722 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	95 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_376_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_376_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_376_Update/ca
      -- 
    ca_849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_376_inst_ack_1, ack => zeropad_CP_182_elements(86)); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	84 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_390_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_390_update_start_
      -- CP-element group 87: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_390_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_390_Sample/ra
      -- CP-element group 87: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_390_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_390_Update/cr
      -- 
    ra_858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_390_inst_ack_0, ack => zeropad_CP_182_elements(87)); -- 
    cr_862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(87), ack => RPIPE_Zeropad_input_pipe_390_inst_req_1); -- 
    -- CP-element group 88:  fork  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: 	91 
    -- CP-element group 88:  members (9) 
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_390_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_390_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_390_Update/ca
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_394_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_394_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_394_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_408_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_408_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_408_Sample/rr
      -- 
    ca_863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_390_inst_ack_1, ack => zeropad_CP_182_elements(88)); -- 
    rr_871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(88), ack => type_cast_394_inst_req_0); -- 
    rr_885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(88), ack => RPIPE_Zeropad_input_pipe_408_inst_req_0); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_394_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_394_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_394_Sample/ra
      -- 
    ra_872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_394_inst_ack_0, ack => zeropad_CP_182_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	722 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	95 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_394_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_394_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_394_Update/ca
      -- 
    ca_877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_394_inst_ack_1, ack => zeropad_CP_182_elements(90)); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	88 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_408_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_408_update_start_
      -- CP-element group 91: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_408_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_408_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_408_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_408_Update/cr
      -- 
    ra_886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_408_inst_ack_0, ack => zeropad_CP_182_elements(91)); -- 
    cr_890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(91), ack => RPIPE_Zeropad_input_pipe_408_inst_req_1); -- 
    -- CP-element group 92:  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (6) 
      -- CP-element group 92: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_408_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_408_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_408_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_412_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_412_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_412_Sample/rr
      -- 
    ca_891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Zeropad_input_pipe_408_inst_ack_1, ack => zeropad_CP_182_elements(92)); -- 
    rr_899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(92), ack => type_cast_412_inst_req_0); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_412_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_412_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_412_Sample/ra
      -- 
    ra_900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_412_inst_ack_0, ack => zeropad_CP_182_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	722 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_412_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_412_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_412_Update/ca
      -- 
    ca_905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_412_inst_ack_1, ack => zeropad_CP_182_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	62 
    -- CP-element group 95: 	66 
    -- CP-element group 95: 	70 
    -- CP-element group 95: 	74 
    -- CP-element group 95: 	78 
    -- CP-element group 95: 	82 
    -- CP-element group 95: 	86 
    -- CP-element group 95: 	90 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Sample/ptr_deref_420_Split/$entry
      -- CP-element group 95: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Sample/ptr_deref_420_Split/$exit
      -- CP-element group 95: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Sample/ptr_deref_420_Split/split_req
      -- CP-element group 95: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Sample/ptr_deref_420_Split/split_ack
      -- CP-element group 95: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Sample/word_access_start/$entry
      -- CP-element group 95: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Sample/word_access_start/word_0/$entry
      -- CP-element group 95: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Sample/word_access_start/word_0/rr
      -- 
    rr_943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(95), ack => ptr_deref_420_store_0_req_0); -- 
    zeropad_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 27) := "zeropad_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(62) & zeropad_CP_182_elements(66) & zeropad_CP_182_elements(70) & zeropad_CP_182_elements(74) & zeropad_CP_182_elements(78) & zeropad_CP_182_elements(82) & zeropad_CP_182_elements(86) & zeropad_CP_182_elements(90) & zeropad_CP_182_elements(94);
      gj_zeropad_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Sample/word_access_start/$exit
      -- CP-element group 96: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Sample/word_access_start/word_0/$exit
      -- CP-element group 96: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Sample/word_access_start/word_0/ra
      -- 
    ra_944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_420_store_0_ack_0, ack => zeropad_CP_182_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	722 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Update/word_access_complete/$exit
      -- CP-element group 97: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Update/word_access_complete/word_0/$exit
      -- CP-element group 97: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Update/word_access_complete/word_0/ca
      -- 
    ca_955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_420_store_0_ack_1, ack => zeropad_CP_182_elements(97)); -- 
    -- CP-element group 98:  branch  join  transition  place  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	59 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (10) 
      -- CP-element group 98: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433__exit__
      -- CP-element group 98: 	 branch_block_stmt_43/if_stmt_434__entry__
      -- CP-element group 98: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/$exit
      -- CP-element group 98: 	 branch_block_stmt_43/if_stmt_434_dead_link/$entry
      -- CP-element group 98: 	 branch_block_stmt_43/if_stmt_434_eval_test/$entry
      -- CP-element group 98: 	 branch_block_stmt_43/if_stmt_434_eval_test/$exit
      -- CP-element group 98: 	 branch_block_stmt_43/if_stmt_434_eval_test/branch_req
      -- CP-element group 98: 	 branch_block_stmt_43/R_exitcond_435_place
      -- CP-element group 98: 	 branch_block_stmt_43/if_stmt_434_if_link/$entry
      -- CP-element group 98: 	 branch_block_stmt_43/if_stmt_434_else_link/$entry
      -- 
    branch_req_963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(98), ack => if_stmt_434_branch_req_0); -- 
    zeropad_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "zeropad_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(59) & zeropad_CP_182_elements(97);
      gj_zeropad_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  merge  transition  place  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	723 
    -- CP-element group 99:  members (13) 
      -- CP-element group 99: 	 branch_block_stmt_43/merge_stmt_440__exit__
      -- CP-element group 99: 	 branch_block_stmt_43/forx_xendx_xloopexit_forx_xend
      -- CP-element group 99: 	 branch_block_stmt_43/if_stmt_434_if_link/$exit
      -- CP-element group 99: 	 branch_block_stmt_43/if_stmt_434_if_link/if_choice_transition
      -- CP-element group 99: 	 branch_block_stmt_43/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 99: 	 branch_block_stmt_43/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 99: 	 branch_block_stmt_43/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 99: 	 branch_block_stmt_43/merge_stmt_440_PhiReqMerge
      -- CP-element group 99: 	 branch_block_stmt_43/merge_stmt_440_PhiAck/$entry
      -- CP-element group 99: 	 branch_block_stmt_43/merge_stmt_440_PhiAck/$exit
      -- CP-element group 99: 	 branch_block_stmt_43/merge_stmt_440_PhiAck/dummy
      -- CP-element group 99: 	 branch_block_stmt_43/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 99: 	 branch_block_stmt_43/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_434_branch_ack_1, ack => zeropad_CP_182_elements(99)); -- 
    -- CP-element group 100:  fork  transition  place  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	718 
    -- CP-element group 100: 	719 
    -- CP-element group 100:  members (12) 
      -- CP-element group 100: 	 branch_block_stmt_43/if_stmt_434_else_link/$exit
      -- CP-element group 100: 	 branch_block_stmt_43/if_stmt_434_else_link/else_choice_transition
      -- CP-element group 100: 	 branch_block_stmt_43/forx_xbody_forx_xbody
      -- CP-element group 100: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 100: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/phi_stmt_269/$entry
      -- CP-element group 100: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_sources/$entry
      -- CP-element group 100: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_275/$entry
      -- CP-element group 100: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_275/SplitProtocol/$entry
      -- CP-element group 100: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_275/SplitProtocol/Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_275/SplitProtocol/Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_275/SplitProtocol/Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_275/SplitProtocol/Update/cr
      -- 
    else_choice_transition_972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_434_branch_ack_0, ack => zeropad_CP_182_elements(100)); -- 
    rr_3339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(100), ack => type_cast_275_inst_req_0); -- 
    cr_3344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(100), ack => type_cast_275_inst_req_1); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	723 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_43/call_stmt_445/call_stmt_445_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_43/call_stmt_445/call_stmt_445_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_43/call_stmt_445/call_stmt_445_Sample/cra
      -- 
    cra_986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_445_call_ack_0, ack => zeropad_CP_182_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	723 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (33) 
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Update/word_access_complete/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Sample/word_access_start/$entry
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Update/word_access_complete/$entry
      -- CP-element group 102: 	 branch_block_stmt_43/call_stmt_445__exit__
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531__entry__
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Sample/word_access_start/word_0/rr
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Sample/word_access_start/word_0/$entry
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_word_addrgen/root_register_ack
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_word_addrgen/root_register_req
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Update/word_access_complete/word_0/cr
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_word_addrgen/$exit
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_word_addrgen/$entry
      -- CP-element group 102: 	 branch_block_stmt_43/call_stmt_445/$exit
      -- CP-element group 102: 	 branch_block_stmt_43/call_stmt_445/call_stmt_445_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_43/call_stmt_445/call_stmt_445_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_43/call_stmt_445/call_stmt_445_Update/cca
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/$entry
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_update_start_
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_base_address_calculated
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_word_address_calculated
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_root_address_calculated
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_base_address_resized
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_base_addr_resize/$entry
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_base_addr_resize/$exit
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_base_addr_resize/base_resize_req
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_base_addr_resize/base_resize_ack
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_base_plus_offset/$entry
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_base_plus_offset/$exit
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_base_plus_offset/sum_rename_req
      -- CP-element group 102: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_base_plus_offset/sum_rename_ack
      -- 
    cca_991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_445_call_ack_1, ack => zeropad_CP_182_elements(102)); -- 
    rr_1027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(102), ack => ptr_deref_491_load_0_req_0); -- 
    cr_1038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(102), ack => ptr_deref_491_load_0_req_1); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (5) 
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Sample/word_access_start/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Sample/word_access_start/word_0/ra
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Sample/word_access_start/word_0/$exit
      -- CP-element group 103: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_sample_completed_
      -- 
    ra_1028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_491_load_0_ack_0, ack => zeropad_CP_182_elements(103)); -- 
    -- CP-element group 104:  fork  transition  place  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	724 
    -- CP-element group 104: 	725 
    -- CP-element group 104: 	727 
    -- CP-element group 104: 	728 
    -- CP-element group 104:  members (29) 
      -- CP-element group 104: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Update/word_access_complete/word_0/$exit
      -- CP-element group 104: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Update/word_access_complete/$exit
      -- CP-element group 104: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531__exit__
      -- CP-element group 104: 	 branch_block_stmt_43/forx_xend_whilex_xbody
      -- CP-element group 104: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Update/ptr_deref_491_Merge/merge_ack
      -- CP-element group 104: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Update/ptr_deref_491_Merge/merge_req
      -- CP-element group 104: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Update/ptr_deref_491_Merge/$exit
      -- CP-element group 104: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Update/ptr_deref_491_Merge/$entry
      -- CP-element group 104: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_Update/word_access_complete/word_0/ca
      -- CP-element group 104: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/$exit
      -- CP-element group 104: 	 branch_block_stmt_43/assign_stmt_451_to_assign_stmt_531/ptr_deref_491_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/$entry
      -- CP-element group 104: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_539/$entry
      -- CP-element group 104: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_539/phi_stmt_539_sources/$entry
      -- CP-element group 104: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_539/phi_stmt_539_sources/type_cast_542/$entry
      -- CP-element group 104: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_539/phi_stmt_539_sources/type_cast_542/SplitProtocol/$entry
      -- CP-element group 104: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_539/phi_stmt_539_sources/type_cast_542/SplitProtocol/Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_539/phi_stmt_539_sources/type_cast_542/SplitProtocol/Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_539/phi_stmt_539_sources/type_cast_542/SplitProtocol/Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_539/phi_stmt_539_sources/type_cast_542/SplitProtocol/Update/cr
      -- CP-element group 104: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_583/$entry
      -- CP-element group 104: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_583/phi_stmt_583_sources/$entry
      -- CP-element group 104: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_586/$entry
      -- CP-element group 104: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_586/SplitProtocol/$entry
      -- CP-element group 104: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_586/SplitProtocol/Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_586/SplitProtocol/Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_586/SplitProtocol/Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_586/SplitProtocol/Update/cr
      -- 
    ca_1039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_491_load_0_ack_1, ack => zeropad_CP_182_elements(104)); -- 
    rr_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(104), ack => type_cast_542_inst_req_0); -- 
    cr_3398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(104), ack => type_cast_542_inst_req_1); -- 
    rr_3416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(104), ack => type_cast_586_inst_req_0); -- 
    cr_3421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(104), ack => type_cast_586_inst_req_1); -- 
    -- CP-element group 105:  transition  place  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	733 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	111 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_43/do_while_stmt_588/$entry
      -- CP-element group 105: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588__entry__
      -- 
    zeropad_CP_182_elements(105) <= zeropad_CP_182_elements(733);
    -- CP-element group 106:  merge  place  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	614 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588__exit__
      -- 
    -- Element group zeropad_CP_182_elements(106) is bound as output of CP function.
    -- CP-element group 107:  merge  place  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_43/do_while_stmt_588/loop_back
      -- 
    -- Element group zeropad_CP_182_elements(107) is bound as output of CP function.
    -- CP-element group 108:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	113 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	612 
    -- CP-element group 108: 	613 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_43/do_while_stmt_588/condition_done
      -- CP-element group 108: 	 branch_block_stmt_43/do_while_stmt_588/loop_exit/$entry
      -- CP-element group 108: 	 branch_block_stmt_43/do_while_stmt_588/loop_taken/$entry
      -- 
    zeropad_CP_182_elements(108) <= zeropad_CP_182_elements(113);
    -- CP-element group 109:  branch  place  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	611 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_43/do_while_stmt_588/loop_body_done
      -- 
    zeropad_CP_182_elements(109) <= zeropad_CP_182_elements(611);
    -- CP-element group 110:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	122 
    -- CP-element group 110: 	143 
    -- CP-element group 110: 	164 
    -- CP-element group 110: 	185 
    -- CP-element group 110: 	206 
    -- CP-element group 110: 	227 
    -- CP-element group 110: 	248 
    -- CP-element group 110: 	269 
    -- CP-element group 110: 	290 
    -- CP-element group 110: 	311 
    -- CP-element group 110: 	332 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/back_edge_to_loop_body
      -- 
    zeropad_CP_182_elements(110) <= zeropad_CP_182_elements(107);
    -- CP-element group 111:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	105 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	124 
    -- CP-element group 111: 	145 
    -- CP-element group 111: 	166 
    -- CP-element group 111: 	187 
    -- CP-element group 111: 	208 
    -- CP-element group 111: 	229 
    -- CP-element group 111: 	250 
    -- CP-element group 111: 	271 
    -- CP-element group 111: 	292 
    -- CP-element group 111: 	313 
    -- CP-element group 111: 	334 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/first_time_through_loop_body
      -- 
    zeropad_CP_182_elements(111) <= zeropad_CP_182_elements(105);
    -- CP-element group 112:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	118 
    -- CP-element group 112: 	119 
    -- CP-element group 112: 	137 
    -- CP-element group 112: 	138 
    -- CP-element group 112: 	158 
    -- CP-element group 112: 	159 
    -- CP-element group 112: 	179 
    -- CP-element group 112: 	180 
    -- CP-element group 112: 	200 
    -- CP-element group 112: 	201 
    -- CP-element group 112: 	221 
    -- CP-element group 112: 	222 
    -- CP-element group 112: 	242 
    -- CP-element group 112: 	243 
    -- CP-element group 112: 	263 
    -- CP-element group 112: 	264 
    -- CP-element group 112: 	284 
    -- CP-element group 112: 	285 
    -- CP-element group 112: 	305 
    -- CP-element group 112: 	306 
    -- CP-element group 112: 	326 
    -- CP-element group 112: 	327 
    -- CP-element group 112: 	388 
    -- CP-element group 112: 	389 
    -- CP-element group 112: 	422 
    -- CP-element group 112: 	563 
    -- CP-element group 112: 	564 
    -- CP-element group 112: 	585 
    -- CP-element group 112: 	609 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/loop_body_start
      -- CP-element group 112: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/$entry
      -- 
    -- Element group zeropad_CP_182_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	117 
    -- CP-element group 113: 	604 
    -- CP-element group 113: 	608 
    -- CP-element group 113: 	609 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	108 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/condition_evaluated
      -- 
    condition_evaluated_1059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(113), ack => do_while_stmt_588_branch_req_0); -- 
    zeropad_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(117) & zeropad_CP_182_elements(604) & zeropad_CP_182_elements(608) & zeropad_CP_182_elements(609);
      gj_zeropad_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	118 
    -- CP-element group 114: 	137 
    -- CP-element group 114: 	158 
    -- CP-element group 114: 	179 
    -- CP-element group 114: 	200 
    -- CP-element group 114: 	221 
    -- CP-element group 114: 	242 
    -- CP-element group 114: 	263 
    -- CP-element group 114: 	284 
    -- CP-element group 114: 	305 
    -- CP-element group 114: 	326 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	117 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	139 
    -- CP-element group 114: 	160 
    -- CP-element group 114: 	181 
    -- CP-element group 114: 	202 
    -- CP-element group 114: 	223 
    -- CP-element group 114: 	244 
    -- CP-element group 114: 	265 
    -- CP-element group 114: 	286 
    -- CP-element group 114: 	307 
    -- CP-element group 114: 	328 
    -- CP-element group 114:  members (2) 
      -- CP-element group 114: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_590_sample_start__ps
      -- CP-element group 114: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/aggregated_phi_sample_req
      -- 
    zeropad_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(118) & zeropad_CP_182_elements(137) & zeropad_CP_182_elements(158) & zeropad_CP_182_elements(179) & zeropad_CP_182_elements(200) & zeropad_CP_182_elements(221) & zeropad_CP_182_elements(242) & zeropad_CP_182_elements(263) & zeropad_CP_182_elements(284) & zeropad_CP_182_elements(305) & zeropad_CP_182_elements(326) & zeropad_CP_182_elements(117);
      gj_zeropad_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	120 
    -- CP-element group 115: 	140 
    -- CP-element group 115: 	161 
    -- CP-element group 115: 	182 
    -- CP-element group 115: 	203 
    -- CP-element group 115: 	224 
    -- CP-element group 115: 	245 
    -- CP-element group 115: 	266 
    -- CP-element group 115: 	287 
    -- CP-element group 115: 	308 
    -- CP-element group 115: 	329 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	364 
    -- CP-element group 115: 	372 
    -- CP-element group 115: 	384 
    -- CP-element group 115: 	399 
    -- CP-element group 115: 	403 
    -- CP-element group 115: 	407 
    -- CP-element group 115: 	443 
    -- CP-element group 115: 	451 
    -- CP-element group 115: 	455 
    -- CP-element group 115: 	463 
    -- CP-element group 115: 	479 
    -- CP-element group 115: 	483 
    -- CP-element group 115: 	487 
    -- CP-element group 115: 	491 
    -- CP-element group 115: 	495 
    -- CP-element group 115: 	499 
    -- CP-element group 115: 	503 
    -- CP-element group 115: 	507 
    -- CP-element group 115: 	515 
    -- CP-element group 115: 	519 
    -- CP-element group 115: 	523 
    -- CP-element group 115: 	527 
    -- CP-element group 115: 	531 
    -- CP-element group 115: 	535 
    -- CP-element group 115: 	539 
    -- CP-element group 115: 	543 
    -- CP-element group 115: 	547 
    -- CP-element group 115: 	551 
    -- CP-element group 115: 	555 
    -- CP-element group 115: 	559 
    -- CP-element group 115: 	574 
    -- CP-element group 115: 	578 
    -- CP-element group 115: 	582 
    -- CP-element group 115: 	586 
    -- CP-element group 115: 	590 
    -- CP-element group 115: 	594 
    -- CP-element group 115: 	598 
    -- CP-element group 115: 	602 
    -- CP-element group 115: 	606 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	118 
    -- CP-element group 115: 	137 
    -- CP-element group 115: 	158 
    -- CP-element group 115: 	179 
    -- CP-element group 115: 	200 
    -- CP-element group 115: 	221 
    -- CP-element group 115: 	242 
    -- CP-element group 115: 	263 
    -- CP-element group 115: 	284 
    -- CP-element group 115: 	305 
    -- CP-element group 115: 	326 
    -- CP-element group 115:  members (12) 
      -- CP-element group 115: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_605_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_595_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_600_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_590_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/aggregated_phi_sample_ack
      -- CP-element group 115: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_610_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_615_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_620_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_625_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_630_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_635_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_640_sample_completed_
      -- 
    zeropad_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(120) & zeropad_CP_182_elements(140) & zeropad_CP_182_elements(161) & zeropad_CP_182_elements(182) & zeropad_CP_182_elements(203) & zeropad_CP_182_elements(224) & zeropad_CP_182_elements(245) & zeropad_CP_182_elements(266) & zeropad_CP_182_elements(287) & zeropad_CP_182_elements(308) & zeropad_CP_182_elements(329);
      gj_zeropad_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	119 
    -- CP-element group 116: 	138 
    -- CP-element group 116: 	159 
    -- CP-element group 116: 	180 
    -- CP-element group 116: 	201 
    -- CP-element group 116: 	222 
    -- CP-element group 116: 	243 
    -- CP-element group 116: 	264 
    -- CP-element group 116: 	285 
    -- CP-element group 116: 	306 
    -- CP-element group 116: 	327 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	141 
    -- CP-element group 116: 	162 
    -- CP-element group 116: 	183 
    -- CP-element group 116: 	204 
    -- CP-element group 116: 	225 
    -- CP-element group 116: 	246 
    -- CP-element group 116: 	267 
    -- CP-element group 116: 	288 
    -- CP-element group 116: 	309 
    -- CP-element group 116: 	330 
    -- CP-element group 116:  members (2) 
      -- CP-element group 116: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_590_update_start__ps
      -- CP-element group 116: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/aggregated_phi_update_req
      -- 
    zeropad_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(119) & zeropad_CP_182_elements(138) & zeropad_CP_182_elements(159) & zeropad_CP_182_elements(180) & zeropad_CP_182_elements(201) & zeropad_CP_182_elements(222) & zeropad_CP_182_elements(243) & zeropad_CP_182_elements(264) & zeropad_CP_182_elements(285) & zeropad_CP_182_elements(306) & zeropad_CP_182_elements(327);
      gj_zeropad_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	121 
    -- CP-element group 117: 	142 
    -- CP-element group 117: 	163 
    -- CP-element group 117: 	184 
    -- CP-element group 117: 	205 
    -- CP-element group 117: 	226 
    -- CP-element group 117: 	247 
    -- CP-element group 117: 	268 
    -- CP-element group 117: 	289 
    -- CP-element group 117: 	310 
    -- CP-element group 117: 	331 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	113 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	114 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/aggregated_phi_update_ack
      -- 
    zeropad_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(121) & zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(184) & zeropad_CP_182_elements(205) & zeropad_CP_182_elements(226) & zeropad_CP_182_elements(247) & zeropad_CP_182_elements(268) & zeropad_CP_182_elements(289) & zeropad_CP_182_elements(310) & zeropad_CP_182_elements(331);
      gj_zeropad_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	112 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	115 
    -- CP-element group 118: 	445 
    -- CP-element group 118: 	453 
    -- CP-element group 118: 	457 
    -- CP-element group 118: 	489 
    -- CP-element group 118: 	537 
    -- CP-element group 118: 	541 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	114 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_590_sample_start_
      -- 
    zeropad_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(115) & zeropad_CP_182_elements(445) & zeropad_CP_182_elements(453) & zeropad_CP_182_elements(457) & zeropad_CP_182_elements(489) & zeropad_CP_182_elements(537) & zeropad_CP_182_elements(541);
      gj_zeropad_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  join  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	112 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	121 
    -- CP-element group 119: 	390 
    -- CP-element group 119: 	536 
    -- CP-element group 119: 	540 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	116 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_590_update_start_
      -- 
    zeropad_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(121) & zeropad_CP_182_elements(390) & zeropad_CP_182_elements(536) & zeropad_CP_182_elements(540);
      gj_zeropad_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	115 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_590_sample_completed__ps
      -- 
    -- Element group zeropad_CP_182_elements(120) is bound as output of CP function.
    -- CP-element group 121:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	117 
    -- CP-element group 121: 	390 
    -- CP-element group 121: 	534 
    -- CP-element group 121: 	538 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	119 
    -- CP-element group 121:  members (15) 
      -- CP-element group 121: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_final_index_sum_regn_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_index_scale_2/scale_rename_req
      -- CP-element group 121: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_index_scale_2/$exit
      -- CP-element group 121: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_index_scale_2/scale_rename_ack
      -- CP-element group 121: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_590_update_completed__ps
      -- CP-element group 121: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_590_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_final_index_sum_regn_Sample/req
      -- CP-element group 121: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_index_scale_2/$entry
      -- CP-element group 121: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_index_resized_2
      -- CP-element group 121: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_index_scaled_2
      -- CP-element group 121: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_index_computed_2
      -- CP-element group 121: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_index_resize_2/$entry
      -- CP-element group 121: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_index_resize_2/$exit
      -- CP-element group 121: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_index_resize_2/index_resize_req
      -- CP-element group 121: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_index_resize_2/index_resize_ack
      -- 
    req_1733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(121), ack => array_obj_ref_789_index_offset_req_0); -- 
    -- Element group zeropad_CP_182_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	110 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_590_loopback_trigger
      -- 
    zeropad_CP_182_elements(122) <= zeropad_CP_182_elements(110);
    -- CP-element group 123:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_590_loopback_sample_req_ps
      -- CP-element group 123: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_590_loopback_sample_req
      -- 
    phi_stmt_590_loopback_sample_req_1074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_590_loopback_sample_req_1074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(123), ack => phi_stmt_590_req_0); -- 
    -- Element group zeropad_CP_182_elements(123) is bound as output of CP function.
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	111 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_590_entry_trigger
      -- 
    zeropad_CP_182_elements(124) <= zeropad_CP_182_elements(111);
    -- CP-element group 125:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_590_entry_sample_req_ps
      -- CP-element group 125: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_590_entry_sample_req
      -- 
    phi_stmt_590_entry_sample_req_1077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_590_entry_sample_req_1077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(125), ack => phi_stmt_590_req_1); -- 
    -- Element group zeropad_CP_182_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_590_phi_mux_ack_ps
      -- CP-element group 126: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_590_phi_mux_ack
      -- 
    phi_stmt_590_phi_mux_ack_1080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_590_ack_0, ack => zeropad_CP_182_elements(126)); -- 
    -- CP-element group 127:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_593_sample_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (1) 
      -- CP-element group 128: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_593_update_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(128) is bound as output of CP function.
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	131 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_593_Sample/rr
      -- CP-element group 129: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_593_Sample/$entry
      -- CP-element group 129: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_593_sample_start_
      -- 
    rr_1093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(129), ack => type_cast_593_inst_req_0); -- 
    zeropad_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(127) & zeropad_CP_182_elements(131);
      gj_zeropad_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	132 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_593_Update/cr
      -- CP-element group 130: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_593_Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_593_update_start_
      -- 
    cr_1098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(130), ack => type_cast_593_inst_req_1); -- 
    zeropad_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(128) & zeropad_CP_182_elements(132);
      gj_zeropad_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	129 
    -- CP-element group 131:  members (4) 
      -- CP-element group 131: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_593_sample_completed__ps
      -- CP-element group 131: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_593_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_593_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_593_sample_completed_
      -- 
    ra_1094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_593_inst_ack_0, ack => zeropad_CP_182_elements(131)); -- 
    -- CP-element group 132:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: marked-successors 
    -- CP-element group 132: 	130 
    -- CP-element group 132:  members (4) 
      -- CP-element group 132: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_593_update_completed__ps
      -- CP-element group 132: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_593_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_593_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_593_update_completed_
      -- 
    ca_1099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_593_inst_ack_1, ack => zeropad_CP_182_elements(132)); -- 
    -- CP-element group 133:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_add_srcx_x1_at_entry_594_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_add_srcx_x1_at_entry_594_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_add_srcx_x1_at_entry_594_sample_completed__ps
      -- CP-element group 133: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_add_srcx_x1_at_entry_594_sample_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(133) is bound as output of CP function.
    -- CP-element group 134:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_add_srcx_x1_at_entry_594_update_start_
      -- CP-element group 134: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_add_srcx_x1_at_entry_594_update_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(134) is bound as output of CP function.
    -- CP-element group 135:  join  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	136 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_add_srcx_x1_at_entry_594_update_completed__ps
      -- 
    zeropad_CP_182_elements(135) <= zeropad_CP_182_elements(136);
    -- CP-element group 136:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	135 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_add_srcx_x1_at_entry_594_update_completed_
      -- 
    -- Element group zeropad_CP_182_elements(136) is a control-delay.
    cp_element_136_delay: control_delay_element  generic map(name => " 136_delay", delay_value => 1)  port map(req => zeropad_CP_182_elements(134), ack => zeropad_CP_182_elements(136), clk => clk, reset =>reset);
    -- CP-element group 137:  join  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	112 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	115 
    -- CP-element group 137: 	465 
    -- CP-element group 137: 	481 
    -- CP-element group 137: 	485 
    -- CP-element group 137: 	493 
    -- CP-element group 137: 	497 
    -- CP-element group 137: 	501 
    -- CP-element group 137: 	505 
    -- CP-element group 137: 	509 
    -- CP-element group 137: 	549 
    -- CP-element group 137: 	553 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	114 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_595_sample_start_
      -- 
    zeropad_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(115) & zeropad_CP_182_elements(465) & zeropad_CP_182_elements(481) & zeropad_CP_182_elements(485) & zeropad_CP_182_elements(493) & zeropad_CP_182_elements(497) & zeropad_CP_182_elements(501) & zeropad_CP_182_elements(505) & zeropad_CP_182_elements(509) & zeropad_CP_182_elements(549) & zeropad_CP_182_elements(553);
      gj_zeropad_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  join  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	112 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	142 
    -- CP-element group 138: 	349 
    -- CP-element group 138: 	353 
    -- CP-element group 138: 	357 
    -- CP-element group 138: 	361 
    -- CP-element group 138: 	369 
    -- CP-element group 138: 	377 
    -- CP-element group 138: 	381 
    -- CP-element group 138: 	396 
    -- CP-element group 138: 	404 
    -- CP-element group 138: 	408 
    -- CP-element group 138: 	412 
    -- CP-element group 138: 	416 
    -- CP-element group 138: 	420 
    -- CP-element group 138: 	428 
    -- CP-element group 138: 	432 
    -- CP-element group 138: 	436 
    -- CP-element group 138: 	468 
    -- CP-element group 138: 	484 
    -- CP-element group 138: 	496 
    -- CP-element group 138: 	504 
    -- CP-element group 138: 	516 
    -- CP-element group 138: 	524 
    -- CP-element group 138: 	528 
    -- CP-element group 138: 	532 
    -- CP-element group 138: 	536 
    -- CP-element group 138: 	540 
    -- CP-element group 138: 	544 
    -- CP-element group 138: 	552 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	116 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_595_update_start_
      -- 
    zeropad_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 29) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1,29 => 1);
      constant place_markings: IntegerArray(0 to 29)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1,29 => 1);
      constant place_delays: IntegerArray(0 to 29) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0,28 => 0,29 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 30); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(142) & zeropad_CP_182_elements(349) & zeropad_CP_182_elements(353) & zeropad_CP_182_elements(357) & zeropad_CP_182_elements(361) & zeropad_CP_182_elements(369) & zeropad_CP_182_elements(377) & zeropad_CP_182_elements(381) & zeropad_CP_182_elements(396) & zeropad_CP_182_elements(404) & zeropad_CP_182_elements(408) & zeropad_CP_182_elements(412) & zeropad_CP_182_elements(416) & zeropad_CP_182_elements(420) & zeropad_CP_182_elements(428) & zeropad_CP_182_elements(432) & zeropad_CP_182_elements(436) & zeropad_CP_182_elements(468) & zeropad_CP_182_elements(484) & zeropad_CP_182_elements(496) & zeropad_CP_182_elements(504) & zeropad_CP_182_elements(516) & zeropad_CP_182_elements(524) & zeropad_CP_182_elements(528) & zeropad_CP_182_elements(532) & zeropad_CP_182_elements(536) & zeropad_CP_182_elements(540) & zeropad_CP_182_elements(544) & zeropad_CP_182_elements(552);
      gj_zeropad_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 30, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	114 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_595_sample_start__ps
      -- 
    zeropad_CP_182_elements(139) <= zeropad_CP_182_elements(114);
    -- CP-element group 140:  join  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	115 
    -- CP-element group 140:  members (1) 
      -- CP-element group 140: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_595_sample_completed__ps
      -- 
    -- Element group zeropad_CP_182_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	116 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_595_update_start__ps
      -- 
    zeropad_CP_182_elements(141) <= zeropad_CP_182_elements(116);
    -- CP-element group 142:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	117 
    -- CP-element group 142: 	347 
    -- CP-element group 142: 	351 
    -- CP-element group 142: 	355 
    -- CP-element group 142: 	359 
    -- CP-element group 142: 	367 
    -- CP-element group 142: 	375 
    -- CP-element group 142: 	379 
    -- CP-element group 142: 	394 
    -- CP-element group 142: 	402 
    -- CP-element group 142: 	406 
    -- CP-element group 142: 	410 
    -- CP-element group 142: 	414 
    -- CP-element group 142: 	418 
    -- CP-element group 142: 	426 
    -- CP-element group 142: 	430 
    -- CP-element group 142: 	434 
    -- CP-element group 142: 	466 
    -- CP-element group 142: 	482 
    -- CP-element group 142: 	494 
    -- CP-element group 142: 	502 
    -- CP-element group 142: 	514 
    -- CP-element group 142: 	522 
    -- CP-element group 142: 	526 
    -- CP-element group 142: 	530 
    -- CP-element group 142: 	534 
    -- CP-element group 142: 	538 
    -- CP-element group 142: 	542 
    -- CP-element group 142: 	550 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	138 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_595_update_completed__ps
      -- CP-element group 142: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_595_update_completed_
      -- 
    -- Element group zeropad_CP_182_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	110 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_595_loopback_trigger
      -- 
    zeropad_CP_182_elements(143) <= zeropad_CP_182_elements(110);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_595_loopback_sample_req_ps
      -- CP-element group 144: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_595_loopback_sample_req
      -- 
    phi_stmt_595_loopback_sample_req_1118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_595_loopback_sample_req_1118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(144), ack => phi_stmt_595_req_0); -- 
    -- Element group zeropad_CP_182_elements(144) is bound as output of CP function.
    -- CP-element group 145:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	111 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (1) 
      -- CP-element group 145: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_595_entry_trigger
      -- 
    zeropad_CP_182_elements(145) <= zeropad_CP_182_elements(111);
    -- CP-element group 146:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (2) 
      -- CP-element group 146: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_595_entry_sample_req_ps
      -- CP-element group 146: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_595_entry_sample_req
      -- 
    phi_stmt_595_entry_sample_req_1121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_595_entry_sample_req_1121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(146), ack => phi_stmt_595_req_1); -- 
    -- Element group zeropad_CP_182_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_595_phi_mux_ack_ps
      -- CP-element group 147: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_595_phi_mux_ack
      -- 
    phi_stmt_595_phi_mux_ack_1124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_595_ack_0, ack => zeropad_CP_182_elements(147)); -- 
    -- CP-element group 148:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_598_sample_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(148) is bound as output of CP function.
    -- CP-element group 149:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_598_update_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(149) is bound as output of CP function.
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_598_Sample/rr
      -- CP-element group 150: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_598_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_598_sample_start_
      -- 
    rr_1137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(150), ack => type_cast_598_inst_req_0); -- 
    zeropad_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(148) & zeropad_CP_182_elements(152);
      gj_zeropad_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_598_Update/cr
      -- CP-element group 151: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_598_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_598_update_start_
      -- 
    cr_1142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(151), ack => type_cast_598_inst_req_1); -- 
    zeropad_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(149) & zeropad_CP_182_elements(153);
      gj_zeropad_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	150 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_598_Sample/ra
      -- CP-element group 152: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_598_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_598_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_598_sample_completed__ps
      -- 
    ra_1138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_598_inst_ack_0, ack => zeropad_CP_182_elements(152)); -- 
    -- CP-element group 153:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	151 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_598_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_598_Update/ca
      -- CP-element group 153: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_598_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_598_update_completed__ps
      -- 
    ca_1143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_598_inst_ack_1, ack => zeropad_CP_182_elements(153)); -- 
    -- CP-element group 154:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (4) 
      -- CP-element group 154: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_target_out_offsetx_x1_at_entry_599_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_target_out_offsetx_x1_at_entry_599_Sample/req
      -- CP-element group 154: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_target_out_offsetx_x1_at_entry_599_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_target_out_offsetx_x1_at_entry_599_sample_start__ps
      -- 
    req_1155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(154), ack => target_out_offsetx_x1_at_entry_539_599_buf_req_0); -- 
    -- Element group zeropad_CP_182_elements(154) is bound as output of CP function.
    -- CP-element group 155:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (4) 
      -- CP-element group 155: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_target_out_offsetx_x1_at_entry_599_Update/req
      -- CP-element group 155: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_target_out_offsetx_x1_at_entry_599_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_target_out_offsetx_x1_at_entry_599_update_start_
      -- CP-element group 155: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_target_out_offsetx_x1_at_entry_599_update_start__ps
      -- 
    req_1160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(155), ack => target_out_offsetx_x1_at_entry_539_599_buf_req_1); -- 
    -- Element group zeropad_CP_182_elements(155) is bound as output of CP function.
    -- CP-element group 156:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (4) 
      -- CP-element group 156: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_target_out_offsetx_x1_at_entry_599_Sample/ack
      -- CP-element group 156: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_target_out_offsetx_x1_at_entry_599_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_target_out_offsetx_x1_at_entry_599_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_target_out_offsetx_x1_at_entry_599_sample_completed__ps
      -- 
    ack_1156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => target_out_offsetx_x1_at_entry_539_599_buf_ack_0, ack => zeropad_CP_182_elements(156)); -- 
    -- CP-element group 157:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157:  members (4) 
      -- CP-element group 157: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_target_out_offsetx_x1_at_entry_599_Update/ack
      -- CP-element group 157: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_target_out_offsetx_x1_at_entry_599_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_target_out_offsetx_x1_at_entry_599_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_target_out_offsetx_x1_at_entry_599_update_completed__ps
      -- 
    ack_1161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => target_out_offsetx_x1_at_entry_539_599_buf_ack_1, ack => zeropad_CP_182_elements(157)); -- 
    -- CP-element group 158:  join  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	112 
    -- CP-element group 158: marked-predecessors 
    -- CP-element group 158: 	115 
    -- CP-element group 158: 	557 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	114 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_600_sample_start_
      -- 
    zeropad_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(115) & zeropad_CP_182_elements(557);
      gj_zeropad_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  join  transition  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	112 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	163 
    -- CP-element group 159: 	349 
    -- CP-element group 159: 	353 
    -- CP-element group 159: 	357 
    -- CP-element group 159: 	361 
    -- CP-element group 159: 	369 
    -- CP-element group 159: 	377 
    -- CP-element group 159: 	381 
    -- CP-element group 159: 	396 
    -- CP-element group 159: 	404 
    -- CP-element group 159: 	408 
    -- CP-element group 159: 	412 
    -- CP-element group 159: 	416 
    -- CP-element group 159: 	420 
    -- CP-element group 159: 	428 
    -- CP-element group 159: 	432 
    -- CP-element group 159: 	436 
    -- CP-element group 159: 	516 
    -- CP-element group 159: 	524 
    -- CP-element group 159: 	528 
    -- CP-element group 159: 	532 
    -- CP-element group 159: 	536 
    -- CP-element group 159: 	540 
    -- CP-element group 159: 	544 
    -- CP-element group 159: 	552 
    -- CP-element group 159: 	556 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	116 
    -- CP-element group 159:  members (1) 
      -- CP-element group 159: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_600_update_start_
      -- 
    zeropad_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 26) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1);
      constant place_markings: IntegerArray(0 to 26)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1);
      constant place_delays: IntegerArray(0 to 26) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 27); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(349) & zeropad_CP_182_elements(353) & zeropad_CP_182_elements(357) & zeropad_CP_182_elements(361) & zeropad_CP_182_elements(369) & zeropad_CP_182_elements(377) & zeropad_CP_182_elements(381) & zeropad_CP_182_elements(396) & zeropad_CP_182_elements(404) & zeropad_CP_182_elements(408) & zeropad_CP_182_elements(412) & zeropad_CP_182_elements(416) & zeropad_CP_182_elements(420) & zeropad_CP_182_elements(428) & zeropad_CP_182_elements(432) & zeropad_CP_182_elements(436) & zeropad_CP_182_elements(516) & zeropad_CP_182_elements(524) & zeropad_CP_182_elements(528) & zeropad_CP_182_elements(532) & zeropad_CP_182_elements(536) & zeropad_CP_182_elements(540) & zeropad_CP_182_elements(544) & zeropad_CP_182_elements(552) & zeropad_CP_182_elements(556);
      gj_zeropad_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 27, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	114 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (1) 
      -- CP-element group 160: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_600_sample_start__ps
      -- 
    zeropad_CP_182_elements(160) <= zeropad_CP_182_elements(114);
    -- CP-element group 161:  join  transition  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	115 
    -- CP-element group 161:  members (1) 
      -- CP-element group 161: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_600_sample_completed__ps
      -- 
    -- Element group zeropad_CP_182_elements(161) is bound as output of CP function.
    -- CP-element group 162:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	116 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (1) 
      -- CP-element group 162: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_600_update_start__ps
      -- 
    zeropad_CP_182_elements(162) <= zeropad_CP_182_elements(116);
    -- CP-element group 163:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	117 
    -- CP-element group 163: 	347 
    -- CP-element group 163: 	351 
    -- CP-element group 163: 	355 
    -- CP-element group 163: 	359 
    -- CP-element group 163: 	367 
    -- CP-element group 163: 	375 
    -- CP-element group 163: 	379 
    -- CP-element group 163: 	394 
    -- CP-element group 163: 	402 
    -- CP-element group 163: 	406 
    -- CP-element group 163: 	410 
    -- CP-element group 163: 	414 
    -- CP-element group 163: 	418 
    -- CP-element group 163: 	426 
    -- CP-element group 163: 	430 
    -- CP-element group 163: 	434 
    -- CP-element group 163: 	514 
    -- CP-element group 163: 	522 
    -- CP-element group 163: 	526 
    -- CP-element group 163: 	530 
    -- CP-element group 163: 	534 
    -- CP-element group 163: 	538 
    -- CP-element group 163: 	542 
    -- CP-element group 163: 	550 
    -- CP-element group 163: 	554 
    -- CP-element group 163: marked-successors 
    -- CP-element group 163: 	159 
    -- CP-element group 163:  members (2) 
      -- CP-element group 163: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_600_update_completed__ps
      -- CP-element group 163: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_600_update_completed_
      -- 
    -- Element group zeropad_CP_182_elements(163) is bound as output of CP function.
    -- CP-element group 164:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	110 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (1) 
      -- CP-element group 164: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_600_loopback_trigger
      -- 
    zeropad_CP_182_elements(164) <= zeropad_CP_182_elements(110);
    -- CP-element group 165:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (2) 
      -- CP-element group 165: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_600_loopback_sample_req_ps
      -- CP-element group 165: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_600_loopback_sample_req
      -- 
    phi_stmt_600_loopback_sample_req_1172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_600_loopback_sample_req_1172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(165), ack => phi_stmt_600_req_0); -- 
    -- Element group zeropad_CP_182_elements(165) is bound as output of CP function.
    -- CP-element group 166:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	111 
    -- CP-element group 166: successors 
    -- CP-element group 166:  members (1) 
      -- CP-element group 166: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_600_entry_trigger
      -- 
    zeropad_CP_182_elements(166) <= zeropad_CP_182_elements(111);
    -- CP-element group 167:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (2) 
      -- CP-element group 167: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_600_entry_sample_req_ps
      -- CP-element group 167: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_600_entry_sample_req
      -- 
    phi_stmt_600_entry_sample_req_1175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_600_entry_sample_req_1175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(167), ack => phi_stmt_600_req_1); -- 
    -- Element group zeropad_CP_182_elements(167) is bound as output of CP function.
    -- CP-element group 168:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (2) 
      -- CP-element group 168: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_600_phi_mux_ack_ps
      -- CP-element group 168: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_600_phi_mux_ack
      -- 
    phi_stmt_600_phi_mux_ack_1178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_600_ack_0, ack => zeropad_CP_182_elements(168)); -- 
    -- CP-element group 169:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (1) 
      -- CP-element group 169: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_603_sample_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(169) is bound as output of CP function.
    -- CP-element group 170:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170:  members (1) 
      -- CP-element group 170: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_603_update_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(170) is bound as output of CP function.
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	173 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_603_Sample/rr
      -- CP-element group 171: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_603_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_603_sample_start_
      -- 
    rr_1191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(171), ack => type_cast_603_inst_req_0); -- 
    zeropad_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(169) & zeropad_CP_182_elements(173);
      gj_zeropad_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	174 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_603_update_start_
      -- CP-element group 172: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_603_Update/cr
      -- CP-element group 172: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_603_Update/$entry
      -- 
    cr_1196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(172), ack => type_cast_603_inst_req_1); -- 
    zeropad_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(170) & zeropad_CP_182_elements(174);
      gj_zeropad_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: marked-successors 
    -- CP-element group 173: 	171 
    -- CP-element group 173:  members (4) 
      -- CP-element group 173: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_603_Sample/ra
      -- CP-element group 173: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_603_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_603_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_603_sample_completed__ps
      -- 
    ra_1192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_603_inst_ack_0, ack => zeropad_CP_182_elements(173)); -- 
    -- CP-element group 174:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: marked-successors 
    -- CP-element group 174: 	172 
    -- CP-element group 174:  members (4) 
      -- CP-element group 174: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_603_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_603_update_completed__ps
      -- CP-element group 174: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_603_Update/ca
      -- CP-element group 174: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_603_Update/$exit
      -- 
    ca_1197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_603_inst_ack_1, ack => zeropad_CP_182_elements(174)); -- 
    -- CP-element group 175:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (4) 
      -- CP-element group 175: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_iNsTr_28_at_entry_604_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_iNsTr_28_at_entry_604_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_iNsTr_28_at_entry_604_sample_completed__ps
      -- CP-element group 175: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_iNsTr_28_at_entry_604_sample_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(175) is bound as output of CP function.
    -- CP-element group 176:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (2) 
      -- CP-element group 176: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_iNsTr_28_at_entry_604_update_start_
      -- CP-element group 176: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_iNsTr_28_at_entry_604_update_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(176) is bound as output of CP function.
    -- CP-element group 177:  join  transition  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	178 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (1) 
      -- CP-element group 177: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_iNsTr_28_at_entry_604_update_completed__ps
      -- 
    zeropad_CP_182_elements(177) <= zeropad_CP_182_elements(178);
    -- CP-element group 178:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	177 
    -- CP-element group 178:  members (1) 
      -- CP-element group 178: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_iNsTr_28_at_entry_604_update_completed_
      -- 
    -- Element group zeropad_CP_182_elements(178) is a control-delay.
    cp_element_178_delay: control_delay_element  generic map(name => " 178_delay", delay_value => 1)  port map(req => zeropad_CP_182_elements(176), ack => zeropad_CP_182_elements(178), clk => clk, reset =>reset);
    -- CP-element group 179:  join  transition  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	112 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	115 
    -- CP-element group 179: 	445 
    -- CP-element group 179: 	453 
    -- CP-element group 179: 	457 
    -- CP-element group 179: 	489 
    -- CP-element group 179: 	517 
    -- CP-element group 179: 	561 
    -- CP-element group 179: 	576 
    -- CP-element group 179: 	580 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	114 
    -- CP-element group 179:  members (1) 
      -- CP-element group 179: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_605_sample_start_
      -- 
    zeropad_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(115) & zeropad_CP_182_elements(445) & zeropad_CP_182_elements(453) & zeropad_CP_182_elements(457) & zeropad_CP_182_elements(489) & zeropad_CP_182_elements(517) & zeropad_CP_182_elements(561) & zeropad_CP_182_elements(576) & zeropad_CP_182_elements(580);
      gj_zeropad_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  join  transition  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	112 
    -- CP-element group 180: marked-predecessors 
    -- CP-element group 180: 	184 
    -- CP-element group 180: 	565 
    -- CP-element group 180: 	575 
    -- CP-element group 180: 	579 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	116 
    -- CP-element group 180:  members (1) 
      -- CP-element group 180: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_605_update_start_
      -- 
    zeropad_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(184) & zeropad_CP_182_elements(565) & zeropad_CP_182_elements(575) & zeropad_CP_182_elements(579);
      gj_zeropad_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	114 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (1) 
      -- CP-element group 181: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_605_sample_start__ps
      -- 
    zeropad_CP_182_elements(181) <= zeropad_CP_182_elements(114);
    -- CP-element group 182:  join  transition  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	115 
    -- CP-element group 182:  members (1) 
      -- CP-element group 182: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_605_sample_completed__ps
      -- 
    -- Element group zeropad_CP_182_elements(182) is bound as output of CP function.
    -- CP-element group 183:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	116 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (1) 
      -- CP-element group 183: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_605_update_start__ps
      -- 
    zeropad_CP_182_elements(183) <= zeropad_CP_182_elements(116);
    -- CP-element group 184:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	117 
    -- CP-element group 184: 	565 
    -- CP-element group 184: 	573 
    -- CP-element group 184: 	577 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	180 
    -- CP-element group 184:  members (15) 
      -- CP-element group 184: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_605_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_605_update_completed__ps
      -- CP-element group 184: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_final_index_sum_regn_Sample/req
      -- CP-element group 184: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_final_index_sum_regn_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_index_scale_2/scale_rename_ack
      -- CP-element group 184: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_index_scale_2/scale_rename_req
      -- CP-element group 184: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_index_scale_2/$exit
      -- CP-element group 184: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_index_scale_2/$entry
      -- CP-element group 184: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_index_resize_2/index_resize_ack
      -- CP-element group 184: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_index_resize_2/index_resize_req
      -- CP-element group 184: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_index_resize_2/$exit
      -- CP-element group 184: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_index_resize_2/$entry
      -- CP-element group 184: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_index_computed_2
      -- CP-element group 184: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_index_scaled_2
      -- CP-element group 184: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_index_resized_2
      -- 
    req_2403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(184), ack => array_obj_ref_1187_index_offset_req_0); -- 
    -- Element group zeropad_CP_182_elements(184) is bound as output of CP function.
    -- CP-element group 185:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	110 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (1) 
      -- CP-element group 185: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_605_loopback_trigger
      -- 
    zeropad_CP_182_elements(185) <= zeropad_CP_182_elements(110);
    -- CP-element group 186:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: successors 
    -- CP-element group 186:  members (2) 
      -- CP-element group 186: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_605_loopback_sample_req_ps
      -- CP-element group 186: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_605_loopback_sample_req
      -- 
    phi_stmt_605_loopback_sample_req_1216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_605_loopback_sample_req_1216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(186), ack => phi_stmt_605_req_0); -- 
    -- Element group zeropad_CP_182_elements(186) is bound as output of CP function.
    -- CP-element group 187:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	111 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (1) 
      -- CP-element group 187: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_605_entry_trigger
      -- 
    zeropad_CP_182_elements(187) <= zeropad_CP_182_elements(111);
    -- CP-element group 188:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (2) 
      -- CP-element group 188: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_605_entry_sample_req_ps
      -- CP-element group 188: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_605_entry_sample_req
      -- 
    phi_stmt_605_entry_sample_req_1219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_605_entry_sample_req_1219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(188), ack => phi_stmt_605_req_1); -- 
    -- Element group zeropad_CP_182_elements(188) is bound as output of CP function.
    -- CP-element group 189:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (2) 
      -- CP-element group 189: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_605_phi_mux_ack_ps
      -- CP-element group 189: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_605_phi_mux_ack
      -- 
    phi_stmt_605_phi_mux_ack_1222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_605_ack_0, ack => zeropad_CP_182_elements(189)); -- 
    -- CP-element group 190:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (1) 
      -- CP-element group 190: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_608_sample_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(190) is bound as output of CP function.
    -- CP-element group 191:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	193 
    -- CP-element group 191:  members (1) 
      -- CP-element group 191: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_608_update_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(191) is bound as output of CP function.
    -- CP-element group 192:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: marked-predecessors 
    -- CP-element group 192: 	194 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	194 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_608_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_608_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_608_Sample/$entry
      -- 
    rr_1235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(192), ack => type_cast_608_inst_req_0); -- 
    zeropad_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(190) & zeropad_CP_182_elements(194);
      gj_zeropad_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	191 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	195 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_608_Update/cr
      -- CP-element group 193: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_608_Update/$entry
      -- CP-element group 193: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_608_update_start_
      -- 
    cr_1240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(193), ack => type_cast_608_inst_req_1); -- 
    zeropad_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(191) & zeropad_CP_182_elements(195);
      gj_zeropad_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	192 
    -- CP-element group 194: successors 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	192 
    -- CP-element group 194:  members (4) 
      -- CP-element group 194: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_608_sample_completed__ps
      -- CP-element group 194: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_608_Sample/ra
      -- CP-element group 194: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_608_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_608_sample_completed_
      -- 
    ra_1236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_608_inst_ack_0, ack => zeropad_CP_182_elements(194)); -- 
    -- CP-element group 195:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	193 
    -- CP-element group 195: successors 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (4) 
      -- CP-element group 195: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_608_update_completed__ps
      -- CP-element group 195: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_608_Update/ca
      -- CP-element group 195: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_608_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_608_update_completed_
      -- 
    ca_1241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_608_inst_ack_1, ack => zeropad_CP_182_elements(195)); -- 
    -- CP-element group 196:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (4) 
      -- CP-element group 196: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_add_outx_x1_at_entry_609_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_add_outx_x1_at_entry_609_sample_completed__ps
      -- CP-element group 196: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_add_outx_x1_at_entry_609_sample_start__ps
      -- CP-element group 196: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_add_outx_x1_at_entry_609_sample_start_
      -- 
    -- Element group zeropad_CP_182_elements(196) is bound as output of CP function.
    -- CP-element group 197:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (2) 
      -- CP-element group 197: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_add_outx_x1_at_entry_609_update_start_
      -- CP-element group 197: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_add_outx_x1_at_entry_609_update_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(197) is bound as output of CP function.
    -- CP-element group 198:  join  transition  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	199 
    -- CP-element group 198: successors 
    -- CP-element group 198:  members (1) 
      -- CP-element group 198: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_add_outx_x1_at_entry_609_update_completed__ps
      -- 
    zeropad_CP_182_elements(198) <= zeropad_CP_182_elements(199);
    -- CP-element group 199:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	198 
    -- CP-element group 199:  members (1) 
      -- CP-element group 199: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_add_outx_x1_at_entry_609_update_completed_
      -- 
    -- Element group zeropad_CP_182_elements(199) is a control-delay.
    cp_element_199_delay: control_delay_element  generic map(name => " 199_delay", delay_value => 1)  port map(req => zeropad_CP_182_elements(197), ack => zeropad_CP_182_elements(199), clk => clk, reset =>reset);
    -- CP-element group 200:  join  transition  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	112 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	115 
    -- CP-element group 200: 	445 
    -- CP-element group 200: 	453 
    -- CP-element group 200: 	457 
    -- CP-element group 200: 	489 
    -- CP-element group 200: 	517 
    -- CP-element group 200: 	561 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	114 
    -- CP-element group 200:  members (1) 
      -- CP-element group 200: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_610_sample_start_
      -- 
    zeropad_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(115) & zeropad_CP_182_elements(445) & zeropad_CP_182_elements(453) & zeropad_CP_182_elements(457) & zeropad_CP_182_elements(489) & zeropad_CP_182_elements(517) & zeropad_CP_182_elements(561);
      gj_zeropad_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  join  transition  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	112 
    -- CP-element group 201: marked-predecessors 
    -- CP-element group 201: 	205 
    -- CP-element group 201: 	560 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	116 
    -- CP-element group 201:  members (1) 
      -- CP-element group 201: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_610_update_start_
      -- 
    zeropad_cp_element_group_201: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_201"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(205) & zeropad_CP_182_elements(560);
      gj_zeropad_cp_element_group_201 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(201), clk => clk, reset => reset); --
    end block;
    -- CP-element group 202:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	114 
    -- CP-element group 202: successors 
    -- CP-element group 202:  members (1) 
      -- CP-element group 202: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_610_sample_start__ps
      -- 
    zeropad_CP_182_elements(202) <= zeropad_CP_182_elements(114);
    -- CP-element group 203:  join  transition  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	115 
    -- CP-element group 203:  members (1) 
      -- CP-element group 203: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_610_sample_completed__ps
      -- 
    -- Element group zeropad_CP_182_elements(203) is bound as output of CP function.
    -- CP-element group 204:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	116 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_610_update_start__ps
      -- 
    zeropad_CP_182_elements(204) <= zeropad_CP_182_elements(116);
    -- CP-element group 205:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	117 
    -- CP-element group 205: 	558 
    -- CP-element group 205: marked-successors 
    -- CP-element group 205: 	201 
    -- CP-element group 205:  members (2) 
      -- CP-element group 205: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_610_update_completed__ps
      -- CP-element group 205: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_610_update_completed_
      -- 
    -- Element group zeropad_CP_182_elements(205) is bound as output of CP function.
    -- CP-element group 206:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	110 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (1) 
      -- CP-element group 206: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_610_loopback_trigger
      -- 
    zeropad_CP_182_elements(206) <= zeropad_CP_182_elements(110);
    -- CP-element group 207:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: successors 
    -- CP-element group 207:  members (2) 
      -- CP-element group 207: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_610_loopback_sample_req_ps
      -- CP-element group 207: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_610_loopback_sample_req
      -- 
    phi_stmt_610_loopback_sample_req_1260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_610_loopback_sample_req_1260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(207), ack => phi_stmt_610_req_0); -- 
    -- Element group zeropad_CP_182_elements(207) is bound as output of CP function.
    -- CP-element group 208:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	111 
    -- CP-element group 208: successors 
    -- CP-element group 208:  members (1) 
      -- CP-element group 208: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_610_entry_trigger
      -- 
    zeropad_CP_182_elements(208) <= zeropad_CP_182_elements(111);
    -- CP-element group 209:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: successors 
    -- CP-element group 209:  members (2) 
      -- CP-element group 209: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_610_entry_sample_req
      -- CP-element group 209: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_610_entry_sample_req_ps
      -- 
    phi_stmt_610_entry_sample_req_1263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_610_entry_sample_req_1263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(209), ack => phi_stmt_610_req_1); -- 
    -- Element group zeropad_CP_182_elements(209) is bound as output of CP function.
    -- CP-element group 210:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: successors 
    -- CP-element group 210:  members (2) 
      -- CP-element group 210: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_610_phi_mux_ack
      -- CP-element group 210: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_610_phi_mux_ack_ps
      -- 
    phi_stmt_610_phi_mux_ack_1266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_610_ack_0, ack => zeropad_CP_182_elements(210)); -- 
    -- CP-element group 211:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (1) 
      -- CP-element group 211: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_613_sample_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(211) is bound as output of CP function.
    -- CP-element group 212:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	214 
    -- CP-element group 212:  members (1) 
      -- CP-element group 212: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_613_update_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(212) is bound as output of CP function.
    -- CP-element group 213:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: marked-predecessors 
    -- CP-element group 213: 	215 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	215 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_613_Sample/rr
      -- CP-element group 213: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_613_Sample/$entry
      -- CP-element group 213: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_613_sample_start_
      -- 
    rr_1279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(213), ack => type_cast_613_inst_req_0); -- 
    zeropad_cp_element_group_213: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_213"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(211) & zeropad_CP_182_elements(215);
      gj_zeropad_cp_element_group_213 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(213), clk => clk, reset => reset); --
    end block;
    -- CP-element group 214:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	212 
    -- CP-element group 214: marked-predecessors 
    -- CP-element group 214: 	216 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_613_update_start_
      -- CP-element group 214: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_613_Update/cr
      -- CP-element group 214: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_613_Update/$entry
      -- 
    cr_1284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(214), ack => type_cast_613_inst_req_1); -- 
    zeropad_cp_element_group_214: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_214"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(212) & zeropad_CP_182_elements(216);
      gj_zeropad_cp_element_group_214 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 215:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	213 
    -- CP-element group 215: successors 
    -- CP-element group 215: marked-successors 
    -- CP-element group 215: 	213 
    -- CP-element group 215:  members (4) 
      -- CP-element group 215: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_613_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_613_sample_completed__ps
      -- CP-element group 215: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_613_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_613_Sample/ra
      -- 
    ra_1280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_613_inst_ack_0, ack => zeropad_CP_182_elements(215)); -- 
    -- CP-element group 216:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: successors 
    -- CP-element group 216: marked-successors 
    -- CP-element group 216: 	214 
    -- CP-element group 216:  members (4) 
      -- CP-element group 216: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_613_update_completed__ps
      -- CP-element group 216: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_613_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_613_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_613_Update/ca
      -- 
    ca_1285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_613_inst_ack_1, ack => zeropad_CP_182_elements(216)); -- 
    -- CP-element group 217:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (4) 
      -- CP-element group 217: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_output_byte_countx_x0_at_entry_614_sample_completed__ps
      -- CP-element group 217: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_output_byte_countx_x0_at_entry_614_sample_start_
      -- CP-element group 217: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_output_byte_countx_x0_at_entry_614_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_output_byte_countx_x0_at_entry_614_sample_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(217) is bound as output of CP function.
    -- CP-element group 218:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218:  members (2) 
      -- CP-element group 218: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_output_byte_countx_x0_at_entry_614_update_start__ps
      -- CP-element group 218: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_output_byte_countx_x0_at_entry_614_update_start_
      -- 
    -- Element group zeropad_CP_182_elements(218) is bound as output of CP function.
    -- CP-element group 219:  join  transition  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	220 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (1) 
      -- CP-element group 219: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_output_byte_countx_x0_at_entry_614_update_completed__ps
      -- 
    zeropad_CP_182_elements(219) <= zeropad_CP_182_elements(220);
    -- CP-element group 220:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	219 
    -- CP-element group 220:  members (1) 
      -- CP-element group 220: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_output_byte_countx_x0_at_entry_614_update_completed_
      -- 
    -- Element group zeropad_CP_182_elements(220) is a control-delay.
    cp_element_220_delay: control_delay_element  generic map(name => " 220_delay", delay_value => 1)  port map(req => zeropad_CP_182_elements(218), ack => zeropad_CP_182_elements(220), clk => clk, reset =>reset);
    -- CP-element group 221:  join  transition  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	112 
    -- CP-element group 221: marked-predecessors 
    -- CP-element group 221: 	115 
    -- CP-element group 221: 	445 
    -- CP-element group 221: 	453 
    -- CP-element group 221: 	457 
    -- CP-element group 221: 	489 
    -- CP-element group 221: 	529 
    -- CP-element group 221: 	533 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	114 
    -- CP-element group 221:  members (1) 
      -- CP-element group 221: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_615_sample_start_
      -- 
    zeropad_cp_element_group_221: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_221"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(115) & zeropad_CP_182_elements(445) & zeropad_CP_182_elements(453) & zeropad_CP_182_elements(457) & zeropad_CP_182_elements(489) & zeropad_CP_182_elements(529) & zeropad_CP_182_elements(533);
      gj_zeropad_cp_element_group_221 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(221), clk => clk, reset => reset); --
    end block;
    -- CP-element group 222:  join  transition  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	112 
    -- CP-element group 222: marked-predecessors 
    -- CP-element group 222: 	226 
    -- CP-element group 222: 	349 
    -- CP-element group 222: 	396 
    -- CP-element group 222: 	404 
    -- CP-element group 222: 	408 
    -- CP-element group 222: 	412 
    -- CP-element group 222: 	416 
    -- CP-element group 222: 	420 
    -- CP-element group 222: 	428 
    -- CP-element group 222: 	432 
    -- CP-element group 222: 	436 
    -- CP-element group 222: 	528 
    -- CP-element group 222: 	532 
    -- CP-element group 222: 	536 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	116 
    -- CP-element group 222:  members (1) 
      -- CP-element group 222: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_615_update_start_
      -- 
    zeropad_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 14) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1);
      constant place_markings: IntegerArray(0 to 14)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1);
      constant place_delays: IntegerArray(0 to 14) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 15); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(226) & zeropad_CP_182_elements(349) & zeropad_CP_182_elements(396) & zeropad_CP_182_elements(404) & zeropad_CP_182_elements(408) & zeropad_CP_182_elements(412) & zeropad_CP_182_elements(416) & zeropad_CP_182_elements(420) & zeropad_CP_182_elements(428) & zeropad_CP_182_elements(432) & zeropad_CP_182_elements(436) & zeropad_CP_182_elements(528) & zeropad_CP_182_elements(532) & zeropad_CP_182_elements(536);
      gj_zeropad_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 15, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	114 
    -- CP-element group 223: successors 
    -- CP-element group 223:  members (1) 
      -- CP-element group 223: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_615_sample_start__ps
      -- 
    zeropad_CP_182_elements(223) <= zeropad_CP_182_elements(114);
    -- CP-element group 224:  join  transition  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	115 
    -- CP-element group 224:  members (1) 
      -- CP-element group 224: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_615_sample_completed__ps
      -- 
    -- Element group zeropad_CP_182_elements(224) is bound as output of CP function.
    -- CP-element group 225:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	116 
    -- CP-element group 225: successors 
    -- CP-element group 225:  members (1) 
      -- CP-element group 225: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_615_update_start__ps
      -- 
    zeropad_CP_182_elements(225) <= zeropad_CP_182_elements(116);
    -- CP-element group 226:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	117 
    -- CP-element group 226: 	347 
    -- CP-element group 226: 	394 
    -- CP-element group 226: 	402 
    -- CP-element group 226: 	406 
    -- CP-element group 226: 	410 
    -- CP-element group 226: 	414 
    -- CP-element group 226: 	418 
    -- CP-element group 226: 	426 
    -- CP-element group 226: 	430 
    -- CP-element group 226: 	434 
    -- CP-element group 226: 	526 
    -- CP-element group 226: 	530 
    -- CP-element group 226: 	534 
    -- CP-element group 226: marked-successors 
    -- CP-element group 226: 	222 
    -- CP-element group 226:  members (2) 
      -- CP-element group 226: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_615_update_completed_
      -- CP-element group 226: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_615_update_completed__ps
      -- 
    -- Element group zeropad_CP_182_elements(226) is bound as output of CP function.
    -- CP-element group 227:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	110 
    -- CP-element group 227: successors 
    -- CP-element group 227:  members (1) 
      -- CP-element group 227: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_615_loopback_trigger
      -- 
    zeropad_CP_182_elements(227) <= zeropad_CP_182_elements(110);
    -- CP-element group 228:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (2) 
      -- CP-element group 228: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_615_loopback_sample_req
      -- CP-element group 228: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_615_loopback_sample_req_ps
      -- 
    phi_stmt_615_loopback_sample_req_1304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_615_loopback_sample_req_1304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(228), ack => phi_stmt_615_req_0); -- 
    -- Element group zeropad_CP_182_elements(228) is bound as output of CP function.
    -- CP-element group 229:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	111 
    -- CP-element group 229: successors 
    -- CP-element group 229:  members (1) 
      -- CP-element group 229: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_615_entry_trigger
      -- 
    zeropad_CP_182_elements(229) <= zeropad_CP_182_elements(111);
    -- CP-element group 230:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: successors 
    -- CP-element group 230:  members (2) 
      -- CP-element group 230: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_615_entry_sample_req
      -- CP-element group 230: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_615_entry_sample_req_ps
      -- 
    phi_stmt_615_entry_sample_req_1307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_615_entry_sample_req_1307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(230), ack => phi_stmt_615_req_1); -- 
    -- Element group zeropad_CP_182_elements(230) is bound as output of CP function.
    -- CP-element group 231:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (2) 
      -- CP-element group 231: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_615_phi_mux_ack
      -- CP-element group 231: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_615_phi_mux_ack_ps
      -- 
    phi_stmt_615_phi_mux_ack_1310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_615_ack_0, ack => zeropad_CP_182_elements(231)); -- 
    -- CP-element group 232:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	234 
    -- CP-element group 232:  members (1) 
      -- CP-element group 232: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_618_sample_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(232) is bound as output of CP function.
    -- CP-element group 233:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (1) 
      -- CP-element group 233: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_618_update_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(233) is bound as output of CP function.
    -- CP-element group 234:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	232 
    -- CP-element group 234: marked-predecessors 
    -- CP-element group 234: 	236 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_618_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_618_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_618_Sample/rr
      -- 
    rr_1323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(234), ack => type_cast_618_inst_req_0); -- 
    zeropad_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(232) & zeropad_CP_182_elements(236);
      gj_zeropad_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: marked-predecessors 
    -- CP-element group 235: 	237 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	237 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_618_update_start_
      -- CP-element group 235: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_618_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_618_Update/cr
      -- 
    cr_1328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(235), ack => type_cast_618_inst_req_1); -- 
    zeropad_cp_element_group_235: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_235"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(233) & zeropad_CP_182_elements(237);
      gj_zeropad_cp_element_group_235 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(235), clk => clk, reset => reset); --
    end block;
    -- CP-element group 236:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236: marked-successors 
    -- CP-element group 236: 	234 
    -- CP-element group 236:  members (4) 
      -- CP-element group 236: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_618_sample_completed__ps
      -- CP-element group 236: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_618_sample_completed_
      -- CP-element group 236: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_618_Sample/$exit
      -- CP-element group 236: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_618_Sample/ra
      -- 
    ra_1324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_618_inst_ack_0, ack => zeropad_CP_182_elements(236)); -- 
    -- CP-element group 237:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	235 
    -- CP-element group 237: successors 
    -- CP-element group 237: marked-successors 
    -- CP-element group 237: 	235 
    -- CP-element group 237:  members (4) 
      -- CP-element group 237: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_618_update_completed__ps
      -- CP-element group 237: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_618_update_completed_
      -- CP-element group 237: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_618_Update/$exit
      -- CP-element group 237: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_618_Update/ca
      -- 
    ca_1329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_618_inst_ack_1, ack => zeropad_CP_182_elements(237)); -- 
    -- CP-element group 238:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: successors 
    -- CP-element group 238:  members (4) 
      -- CP-element group 238: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_byte_countx_x1_at_entry_619_sample_start__ps
      -- CP-element group 238: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_byte_countx_x1_at_entry_619_sample_completed__ps
      -- CP-element group 238: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_byte_countx_x1_at_entry_619_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_byte_countx_x1_at_entry_619_sample_completed_
      -- 
    -- Element group zeropad_CP_182_elements(238) is bound as output of CP function.
    -- CP-element group 239:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	241 
    -- CP-element group 239:  members (2) 
      -- CP-element group 239: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_byte_countx_x1_at_entry_619_update_start__ps
      -- CP-element group 239: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_byte_countx_x1_at_entry_619_update_start_
      -- 
    -- Element group zeropad_CP_182_elements(239) is bound as output of CP function.
    -- CP-element group 240:  join  transition  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	241 
    -- CP-element group 240: successors 
    -- CP-element group 240:  members (1) 
      -- CP-element group 240: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_byte_countx_x1_at_entry_619_update_completed__ps
      -- 
    zeropad_CP_182_elements(240) <= zeropad_CP_182_elements(241);
    -- CP-element group 241:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	239 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	240 
    -- CP-element group 241:  members (1) 
      -- CP-element group 241: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_byte_countx_x1_at_entry_619_update_completed_
      -- 
    -- Element group zeropad_CP_182_elements(241) is a control-delay.
    cp_element_241_delay: control_delay_element  generic map(name => " 241_delay", delay_value => 1)  port map(req => zeropad_CP_182_elements(239), ack => zeropad_CP_182_elements(241), clk => clk, reset =>reset);
    -- CP-element group 242:  join  transition  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	112 
    -- CP-element group 242: marked-predecessors 
    -- CP-element group 242: 	115 
    -- CP-element group 242: 	604 
    -- CP-element group 242: 	608 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	114 
    -- CP-element group 242:  members (1) 
      -- CP-element group 242: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_620_sample_start_
      -- 
    zeropad_cp_element_group_242: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_242"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(115) & zeropad_CP_182_elements(604) & zeropad_CP_182_elements(608);
      gj_zeropad_cp_element_group_242 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(242), clk => clk, reset => reset); --
    end block;
    -- CP-element group 243:  join  transition  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	112 
    -- CP-element group 243: marked-predecessors 
    -- CP-element group 243: 	247 
    -- CP-element group 243: 	412 
    -- CP-element group 243: 	607 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	116 
    -- CP-element group 243:  members (1) 
      -- CP-element group 243: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_620_update_start_
      -- 
    zeropad_cp_element_group_243: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_243"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(247) & zeropad_CP_182_elements(412) & zeropad_CP_182_elements(607);
      gj_zeropad_cp_element_group_243 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(243), clk => clk, reset => reset); --
    end block;
    -- CP-element group 244:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	114 
    -- CP-element group 244: successors 
    -- CP-element group 244:  members (1) 
      -- CP-element group 244: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_620_sample_start__ps
      -- 
    zeropad_CP_182_elements(244) <= zeropad_CP_182_elements(114);
    -- CP-element group 245:  join  transition  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	115 
    -- CP-element group 245:  members (1) 
      -- CP-element group 245: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_620_sample_completed__ps
      -- 
    -- Element group zeropad_CP_182_elements(245) is bound as output of CP function.
    -- CP-element group 246:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	116 
    -- CP-element group 246: successors 
    -- CP-element group 246:  members (1) 
      -- CP-element group 246: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_620_update_start__ps
      -- 
    zeropad_CP_182_elements(246) <= zeropad_CP_182_elements(116);
    -- CP-element group 247:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	117 
    -- CP-element group 247: 	410 
    -- CP-element group 247: 	605 
    -- CP-element group 247: marked-successors 
    -- CP-element group 247: 	243 
    -- CP-element group 247:  members (2) 
      -- CP-element group 247: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_620_update_completed_
      -- CP-element group 247: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_620_update_completed__ps
      -- 
    -- Element group zeropad_CP_182_elements(247) is bound as output of CP function.
    -- CP-element group 248:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	110 
    -- CP-element group 248: successors 
    -- CP-element group 248:  members (1) 
      -- CP-element group 248: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_620_loopback_trigger
      -- 
    zeropad_CP_182_elements(248) <= zeropad_CP_182_elements(110);
    -- CP-element group 249:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: successors 
    -- CP-element group 249:  members (2) 
      -- CP-element group 249: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_620_loopback_sample_req
      -- CP-element group 249: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_620_loopback_sample_req_ps
      -- 
    phi_stmt_620_loopback_sample_req_1348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_620_loopback_sample_req_1348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(249), ack => phi_stmt_620_req_0); -- 
    -- Element group zeropad_CP_182_elements(249) is bound as output of CP function.
    -- CP-element group 250:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	111 
    -- CP-element group 250: successors 
    -- CP-element group 250:  members (1) 
      -- CP-element group 250: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_620_entry_trigger
      -- 
    zeropad_CP_182_elements(250) <= zeropad_CP_182_elements(111);
    -- CP-element group 251:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: successors 
    -- CP-element group 251:  members (2) 
      -- CP-element group 251: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_620_entry_sample_req
      -- CP-element group 251: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_620_entry_sample_req_ps
      -- 
    phi_stmt_620_entry_sample_req_1351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_620_entry_sample_req_1351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(251), ack => phi_stmt_620_req_1); -- 
    -- Element group zeropad_CP_182_elements(251) is bound as output of CP function.
    -- CP-element group 252:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: successors 
    -- CP-element group 252:  members (2) 
      -- CP-element group 252: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_620_phi_mux_ack
      -- CP-element group 252: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_620_phi_mux_ack_ps
      -- 
    phi_stmt_620_phi_mux_ack_1354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_620_ack_0, ack => zeropad_CP_182_elements(252)); -- 
    -- CP-element group 253:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (1) 
      -- CP-element group 253: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_623_sample_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(253) is bound as output of CP function.
    -- CP-element group 254:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254:  members (1) 
      -- CP-element group 254: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_623_update_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(254) is bound as output of CP function.
    -- CP-element group 255:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: marked-predecessors 
    -- CP-element group 255: 	257 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	257 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_623_sample_start_
      -- CP-element group 255: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_623_Sample/$entry
      -- CP-element group 255: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_623_Sample/rr
      -- 
    rr_1367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(255), ack => type_cast_623_inst_req_0); -- 
    zeropad_cp_element_group_255: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_255"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(253) & zeropad_CP_182_elements(257);
      gj_zeropad_cp_element_group_255 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(255), clk => clk, reset => reset); --
    end block;
    -- CP-element group 256:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: marked-predecessors 
    -- CP-element group 256: 	258 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	258 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_623_update_start_
      -- CP-element group 256: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_623_Update/$entry
      -- CP-element group 256: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_623_Update/cr
      -- 
    cr_1372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(256), ack => type_cast_623_inst_req_1); -- 
    zeropad_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(254) & zeropad_CP_182_elements(258);
      gj_zeropad_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	255 
    -- CP-element group 257: successors 
    -- CP-element group 257: marked-successors 
    -- CP-element group 257: 	255 
    -- CP-element group 257:  members (4) 
      -- CP-element group 257: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_623_sample_completed__ps
      -- CP-element group 257: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_623_sample_completed_
      -- CP-element group 257: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_623_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_623_Sample/ra
      -- 
    ra_1368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_623_inst_ack_0, ack => zeropad_CP_182_elements(257)); -- 
    -- CP-element group 258:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	256 
    -- CP-element group 258: successors 
    -- CP-element group 258: marked-successors 
    -- CP-element group 258: 	256 
    -- CP-element group 258:  members (4) 
      -- CP-element group 258: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_623_update_completed__ps
      -- CP-element group 258: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_623_update_completed_
      -- CP-element group 258: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_623_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_623_Update/ca
      -- 
    ca_1373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_623_inst_ack_1, ack => zeropad_CP_182_elements(258)); -- 
    -- CP-element group 259:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: successors 
    -- CP-element group 259:  members (4) 
      -- CP-element group 259: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o0x_x1_at_entry_624_sample_start__ps
      -- CP-element group 259: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o0x_x1_at_entry_624_sample_completed__ps
      -- CP-element group 259: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o0x_x1_at_entry_624_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o0x_x1_at_entry_624_sample_completed_
      -- 
    -- Element group zeropad_CP_182_elements(259) is bound as output of CP function.
    -- CP-element group 260:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	262 
    -- CP-element group 260:  members (2) 
      -- CP-element group 260: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o0x_x1_at_entry_624_update_start__ps
      -- CP-element group 260: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o0x_x1_at_entry_624_update_start_
      -- 
    -- Element group zeropad_CP_182_elements(260) is bound as output of CP function.
    -- CP-element group 261:  join  transition  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	262 
    -- CP-element group 261: successors 
    -- CP-element group 261:  members (1) 
      -- CP-element group 261: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o0x_x1_at_entry_624_update_completed__ps
      -- 
    zeropad_CP_182_elements(261) <= zeropad_CP_182_elements(262);
    -- CP-element group 262:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	260 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	261 
    -- CP-element group 262:  members (1) 
      -- CP-element group 262: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o0x_x1_at_entry_624_update_completed_
      -- 
    -- Element group zeropad_CP_182_elements(262) is a control-delay.
    cp_element_262_delay: control_delay_element  generic map(name => " 262_delay", delay_value => 1)  port map(req => zeropad_CP_182_elements(260), ack => zeropad_CP_182_elements(262), clk => clk, reset =>reset);
    -- CP-element group 263:  join  transition  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	112 
    -- CP-element group 263: marked-predecessors 
    -- CP-element group 263: 	115 
    -- CP-element group 263: 	592 
    -- CP-element group 263: 	596 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	114 
    -- CP-element group 263:  members (1) 
      -- CP-element group 263: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_625_sample_start_
      -- 
    zeropad_cp_element_group_263: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_263"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(115) & zeropad_CP_182_elements(592) & zeropad_CP_182_elements(596);
      gj_zeropad_cp_element_group_263 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(263), clk => clk, reset => reset); --
    end block;
    -- CP-element group 264:  join  transition  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	112 
    -- CP-element group 264: marked-predecessors 
    -- CP-element group 264: 	268 
    -- CP-element group 264: 	440 
    -- CP-element group 264: 	595 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	116 
    -- CP-element group 264:  members (1) 
      -- CP-element group 264: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_625_update_start_
      -- 
    zeropad_cp_element_group_264: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_264"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(268) & zeropad_CP_182_elements(440) & zeropad_CP_182_elements(595);
      gj_zeropad_cp_element_group_264 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(264), clk => clk, reset => reset); --
    end block;
    -- CP-element group 265:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	114 
    -- CP-element group 265: successors 
    -- CP-element group 265:  members (1) 
      -- CP-element group 265: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_625_sample_start__ps
      -- 
    zeropad_CP_182_elements(265) <= zeropad_CP_182_elements(114);
    -- CP-element group 266:  join  transition  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	115 
    -- CP-element group 266:  members (1) 
      -- CP-element group 266: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_625_sample_completed__ps
      -- 
    -- Element group zeropad_CP_182_elements(266) is bound as output of CP function.
    -- CP-element group 267:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	116 
    -- CP-element group 267: successors 
    -- CP-element group 267:  members (1) 
      -- CP-element group 267: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_625_update_start__ps
      -- 
    zeropad_CP_182_elements(267) <= zeropad_CP_182_elements(116);
    -- CP-element group 268:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	117 
    -- CP-element group 268: 	438 
    -- CP-element group 268: 	593 
    -- CP-element group 268: marked-successors 
    -- CP-element group 268: 	264 
    -- CP-element group 268:  members (2) 
      -- CP-element group 268: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_625_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_625_update_completed__ps
      -- 
    -- Element group zeropad_CP_182_elements(268) is bound as output of CP function.
    -- CP-element group 269:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	110 
    -- CP-element group 269: successors 
    -- CP-element group 269:  members (1) 
      -- CP-element group 269: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_625_loopback_trigger
      -- 
    zeropad_CP_182_elements(269) <= zeropad_CP_182_elements(110);
    -- CP-element group 270:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: successors 
    -- CP-element group 270:  members (2) 
      -- CP-element group 270: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_625_loopback_sample_req
      -- CP-element group 270: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_625_loopback_sample_req_ps
      -- 
    phi_stmt_625_loopback_sample_req_1392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_625_loopback_sample_req_1392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(270), ack => phi_stmt_625_req_0); -- 
    -- Element group zeropad_CP_182_elements(270) is bound as output of CP function.
    -- CP-element group 271:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	111 
    -- CP-element group 271: successors 
    -- CP-element group 271:  members (1) 
      -- CP-element group 271: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_625_entry_trigger
      -- 
    zeropad_CP_182_elements(271) <= zeropad_CP_182_elements(111);
    -- CP-element group 272:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: successors 
    -- CP-element group 272:  members (2) 
      -- CP-element group 272: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_625_entry_sample_req
      -- CP-element group 272: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_625_entry_sample_req_ps
      -- 
    phi_stmt_625_entry_sample_req_1395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_625_entry_sample_req_1395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(272), ack => phi_stmt_625_req_1); -- 
    -- Element group zeropad_CP_182_elements(272) is bound as output of CP function.
    -- CP-element group 273:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: successors 
    -- CP-element group 273:  members (2) 
      -- CP-element group 273: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_625_phi_mux_ack
      -- CP-element group 273: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_625_phi_mux_ack_ps
      -- 
    phi_stmt_625_phi_mux_ack_1398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_625_ack_0, ack => zeropad_CP_182_elements(273)); -- 
    -- CP-element group 274:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	276 
    -- CP-element group 274:  members (1) 
      -- CP-element group 274: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_628_sample_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(274) is bound as output of CP function.
    -- CP-element group 275:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	277 
    -- CP-element group 275:  members (1) 
      -- CP-element group 275: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_628_update_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(275) is bound as output of CP function.
    -- CP-element group 276:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: marked-predecessors 
    -- CP-element group 276: 	278 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	278 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_628_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_628_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_628_Sample/rr
      -- 
    rr_1411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(276), ack => type_cast_628_inst_req_0); -- 
    zeropad_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(274) & zeropad_CP_182_elements(278);
      gj_zeropad_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	275 
    -- CP-element group 277: marked-predecessors 
    -- CP-element group 277: 	279 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_628_update_start_
      -- CP-element group 277: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_628_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_628_Update/cr
      -- 
    cr_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(277), ack => type_cast_628_inst_req_1); -- 
    zeropad_cp_element_group_277: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_277"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(275) & zeropad_CP_182_elements(279);
      gj_zeropad_cp_element_group_277 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 278:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	276 
    -- CP-element group 278: successors 
    -- CP-element group 278: marked-successors 
    -- CP-element group 278: 	276 
    -- CP-element group 278:  members (4) 
      -- CP-element group 278: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_628_sample_completed__ps
      -- CP-element group 278: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_628_sample_completed_
      -- CP-element group 278: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_628_Sample/$exit
      -- CP-element group 278: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_628_Sample/ra
      -- 
    ra_1412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_628_inst_ack_0, ack => zeropad_CP_182_elements(278)); -- 
    -- CP-element group 279:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: successors 
    -- CP-element group 279: marked-successors 
    -- CP-element group 279: 	277 
    -- CP-element group 279:  members (4) 
      -- CP-element group 279: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_628_update_completed__ps
      -- CP-element group 279: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_628_update_completed_
      -- CP-element group 279: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_628_Update/$exit
      -- CP-element group 279: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_628_Update/ca
      -- 
    ca_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_628_inst_ack_1, ack => zeropad_CP_182_elements(279)); -- 
    -- CP-element group 280:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: successors 
    -- CP-element group 280:  members (4) 
      -- CP-element group 280: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o1x_x1_at_entry_629_sample_start__ps
      -- CP-element group 280: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o1x_x1_at_entry_629_sample_completed__ps
      -- CP-element group 280: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o1x_x1_at_entry_629_sample_start_
      -- CP-element group 280: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o1x_x1_at_entry_629_sample_completed_
      -- 
    -- Element group zeropad_CP_182_elements(280) is bound as output of CP function.
    -- CP-element group 281:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	283 
    -- CP-element group 281:  members (2) 
      -- CP-element group 281: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o1x_x1_at_entry_629_update_start__ps
      -- CP-element group 281: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o1x_x1_at_entry_629_update_start_
      -- 
    -- Element group zeropad_CP_182_elements(281) is bound as output of CP function.
    -- CP-element group 282:  join  transition  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	283 
    -- CP-element group 282: successors 
    -- CP-element group 282:  members (1) 
      -- CP-element group 282: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o1x_x1_at_entry_629_update_completed__ps
      -- 
    zeropad_CP_182_elements(282) <= zeropad_CP_182_elements(283);
    -- CP-element group 283:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	281 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	282 
    -- CP-element group 283:  members (1) 
      -- CP-element group 283: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o1x_x1_at_entry_629_update_completed_
      -- 
    -- Element group zeropad_CP_182_elements(283) is a control-delay.
    cp_element_283_delay: control_delay_element  generic map(name => " 283_delay", delay_value => 1)  port map(req => zeropad_CP_182_elements(281), ack => zeropad_CP_182_elements(283), clk => clk, reset =>reset);
    -- CP-element group 284:  join  transition  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	112 
    -- CP-element group 284: marked-predecessors 
    -- CP-element group 284: 	115 
    -- CP-element group 284: 	584 
    -- CP-element group 284: 	588 
    -- CP-element group 284: 	600 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	114 
    -- CP-element group 284:  members (1) 
      -- CP-element group 284: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_630_sample_start_
      -- 
    zeropad_cp_element_group_284: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_284"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(115) & zeropad_CP_182_elements(584) & zeropad_CP_182_elements(588) & zeropad_CP_182_elements(600);
      gj_zeropad_cp_element_group_284 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(284), clk => clk, reset => reset); --
    end block;
    -- CP-element group 285:  join  transition  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	112 
    -- CP-element group 285: marked-predecessors 
    -- CP-element group 285: 	289 
    -- CP-element group 285: 	460 
    -- CP-element group 285: 	583 
    -- CP-element group 285: 	599 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	116 
    -- CP-element group 285:  members (1) 
      -- CP-element group 285: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_630_update_start_
      -- 
    zeropad_cp_element_group_285: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_285"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(289) & zeropad_CP_182_elements(460) & zeropad_CP_182_elements(583) & zeropad_CP_182_elements(599);
      gj_zeropad_cp_element_group_285 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(285), clk => clk, reset => reset); --
    end block;
    -- CP-element group 286:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	114 
    -- CP-element group 286: successors 
    -- CP-element group 286:  members (1) 
      -- CP-element group 286: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_630_sample_start__ps
      -- 
    zeropad_CP_182_elements(286) <= zeropad_CP_182_elements(114);
    -- CP-element group 287:  join  transition  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	115 
    -- CP-element group 287:  members (1) 
      -- CP-element group 287: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_630_sample_completed__ps
      -- 
    -- Element group zeropad_CP_182_elements(287) is bound as output of CP function.
    -- CP-element group 288:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	116 
    -- CP-element group 288: successors 
    -- CP-element group 288:  members (1) 
      -- CP-element group 288: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_630_update_start__ps
      -- 
    zeropad_CP_182_elements(288) <= zeropad_CP_182_elements(116);
    -- CP-element group 289:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	117 
    -- CP-element group 289: 	458 
    -- CP-element group 289: 	581 
    -- CP-element group 289: 	597 
    -- CP-element group 289: marked-successors 
    -- CP-element group 289: 	285 
    -- CP-element group 289:  members (2) 
      -- CP-element group 289: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_630_update_completed_
      -- CP-element group 289: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_630_update_completed__ps
      -- 
    -- Element group zeropad_CP_182_elements(289) is bound as output of CP function.
    -- CP-element group 290:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	110 
    -- CP-element group 290: successors 
    -- CP-element group 290:  members (1) 
      -- CP-element group 290: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_630_loopback_trigger
      -- 
    zeropad_CP_182_elements(290) <= zeropad_CP_182_elements(110);
    -- CP-element group 291:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: successors 
    -- CP-element group 291:  members (2) 
      -- CP-element group 291: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_630_loopback_sample_req
      -- CP-element group 291: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_630_loopback_sample_req_ps
      -- 
    phi_stmt_630_loopback_sample_req_1436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_630_loopback_sample_req_1436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(291), ack => phi_stmt_630_req_0); -- 
    -- Element group zeropad_CP_182_elements(291) is bound as output of CP function.
    -- CP-element group 292:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	111 
    -- CP-element group 292: successors 
    -- CP-element group 292:  members (1) 
      -- CP-element group 292: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_630_entry_trigger
      -- 
    zeropad_CP_182_elements(292) <= zeropad_CP_182_elements(111);
    -- CP-element group 293:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: successors 
    -- CP-element group 293:  members (2) 
      -- CP-element group 293: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_630_entry_sample_req
      -- CP-element group 293: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_630_entry_sample_req_ps
      -- 
    phi_stmt_630_entry_sample_req_1439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_630_entry_sample_req_1439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(293), ack => phi_stmt_630_req_1); -- 
    -- Element group zeropad_CP_182_elements(293) is bound as output of CP function.
    -- CP-element group 294:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: successors 
    -- CP-element group 294:  members (2) 
      -- CP-element group 294: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_630_phi_mux_ack
      -- CP-element group 294: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_630_phi_mux_ack_ps
      -- 
    phi_stmt_630_phi_mux_ack_1442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_630_ack_0, ack => zeropad_CP_182_elements(294)); -- 
    -- CP-element group 295:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	297 
    -- CP-element group 295:  members (1) 
      -- CP-element group 295: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_633_sample_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(295) is bound as output of CP function.
    -- CP-element group 296:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	298 
    -- CP-element group 296:  members (1) 
      -- CP-element group 296: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_633_update_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(296) is bound as output of CP function.
    -- CP-element group 297:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	295 
    -- CP-element group 297: marked-predecessors 
    -- CP-element group 297: 	299 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	299 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_633_sample_start_
      -- CP-element group 297: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_633_Sample/$entry
      -- CP-element group 297: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_633_Sample/rr
      -- 
    rr_1455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(297), ack => type_cast_633_inst_req_0); -- 
    zeropad_cp_element_group_297: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_297"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(295) & zeropad_CP_182_elements(299);
      gj_zeropad_cp_element_group_297 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(297), clk => clk, reset => reset); --
    end block;
    -- CP-element group 298:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	296 
    -- CP-element group 298: marked-predecessors 
    -- CP-element group 298: 	300 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	300 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_633_update_start_
      -- CP-element group 298: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_633_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_633_Update/cr
      -- 
    cr_1460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(298), ack => type_cast_633_inst_req_1); -- 
    zeropad_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(296) & zeropad_CP_182_elements(300);
      gj_zeropad_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	297 
    -- CP-element group 299: successors 
    -- CP-element group 299: marked-successors 
    -- CP-element group 299: 	297 
    -- CP-element group 299:  members (4) 
      -- CP-element group 299: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_633_sample_completed__ps
      -- CP-element group 299: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_633_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_633_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_633_Sample/ra
      -- 
    ra_1456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_633_inst_ack_0, ack => zeropad_CP_182_elements(299)); -- 
    -- CP-element group 300:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	298 
    -- CP-element group 300: successors 
    -- CP-element group 300: marked-successors 
    -- CP-element group 300: 	298 
    -- CP-element group 300:  members (4) 
      -- CP-element group 300: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_633_update_completed__ps
      -- CP-element group 300: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_633_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_633_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_633_Update/ca
      -- 
    ca_1461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_633_inst_ack_1, ack => zeropad_CP_182_elements(300)); -- 
    -- CP-element group 301:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: successors 
    -- CP-element group 301:  members (4) 
      -- CP-element group 301: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o2x_x1_at_entry_634_sample_start__ps
      -- CP-element group 301: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o2x_x1_at_entry_634_sample_completed__ps
      -- CP-element group 301: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o2x_x1_at_entry_634_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o2x_x1_at_entry_634_sample_completed_
      -- 
    -- Element group zeropad_CP_182_elements(301) is bound as output of CP function.
    -- CP-element group 302:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	304 
    -- CP-element group 302:  members (2) 
      -- CP-element group 302: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o2x_x1_at_entry_634_update_start__ps
      -- CP-element group 302: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o2x_x1_at_entry_634_update_start_
      -- 
    -- Element group zeropad_CP_182_elements(302) is bound as output of CP function.
    -- CP-element group 303:  join  transition  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	304 
    -- CP-element group 303: successors 
    -- CP-element group 303:  members (1) 
      -- CP-element group 303: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o2x_x1_at_entry_634_update_completed__ps
      -- 
    zeropad_CP_182_elements(303) <= zeropad_CP_182_elements(304);
    -- CP-element group 304:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	302 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	303 
    -- CP-element group 304:  members (1) 
      -- CP-element group 304: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_o2x_x1_at_entry_634_update_completed_
      -- 
    -- Element group zeropad_CP_182_elements(304) is a control-delay.
    cp_element_304_delay: control_delay_element  generic map(name => " 304_delay", delay_value => 1)  port map(req => zeropad_CP_182_elements(302), ack => zeropad_CP_182_elements(304), clk => clk, reset =>reset);
    -- CP-element group 305:  join  transition  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	112 
    -- CP-element group 305: marked-predecessors 
    -- CP-element group 305: 	115 
    -- CP-element group 305: 	366 
    -- CP-element group 305: 	374 
    -- CP-element group 305: 	386 
    -- CP-element group 305: 	445 
    -- CP-element group 305: 	453 
    -- CP-element group 305: 	457 
    -- CP-element group 305: 	489 
    -- CP-element group 305: 	517 
    -- CP-element group 305: 	545 
    -- CP-element group 305: 	561 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	114 
    -- CP-element group 305:  members (1) 
      -- CP-element group 305: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_635_sample_start_
      -- 
    zeropad_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(115) & zeropad_CP_182_elements(366) & zeropad_CP_182_elements(374) & zeropad_CP_182_elements(386) & zeropad_CP_182_elements(445) & zeropad_CP_182_elements(453) & zeropad_CP_182_elements(457) & zeropad_CP_182_elements(489) & zeropad_CP_182_elements(517) & zeropad_CP_182_elements(545) & zeropad_CP_182_elements(561);
      gj_zeropad_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  join  transition  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	112 
    -- CP-element group 306: marked-predecessors 
    -- CP-element group 306: 	310 
    -- CP-element group 306: 	385 
    -- CP-element group 306: 	544 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	116 
    -- CP-element group 306:  members (1) 
      -- CP-element group 306: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_635_update_start_
      -- 
    zeropad_cp_element_group_306: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_306"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(310) & zeropad_CP_182_elements(385) & zeropad_CP_182_elements(544);
      gj_zeropad_cp_element_group_306 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(306), clk => clk, reset => reset); --
    end block;
    -- CP-element group 307:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	114 
    -- CP-element group 307: successors 
    -- CP-element group 307:  members (1) 
      -- CP-element group 307: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_635_sample_start__ps
      -- 
    zeropad_CP_182_elements(307) <= zeropad_CP_182_elements(114);
    -- CP-element group 308:  join  transition  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	115 
    -- CP-element group 308:  members (1) 
      -- CP-element group 308: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_635_sample_completed__ps
      -- 
    -- Element group zeropad_CP_182_elements(308) is bound as output of CP function.
    -- CP-element group 309:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	116 
    -- CP-element group 309: successors 
    -- CP-element group 309:  members (1) 
      -- CP-element group 309: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_635_update_start__ps
      -- 
    zeropad_CP_182_elements(309) <= zeropad_CP_182_elements(116);
    -- CP-element group 310:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	117 
    -- CP-element group 310: 	383 
    -- CP-element group 310: 	542 
    -- CP-element group 310: marked-successors 
    -- CP-element group 310: 	306 
    -- CP-element group 310:  members (2) 
      -- CP-element group 310: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_635_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_635_update_completed__ps
      -- 
    -- Element group zeropad_CP_182_elements(310) is bound as output of CP function.
    -- CP-element group 311:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	110 
    -- CP-element group 311: successors 
    -- CP-element group 311:  members (1) 
      -- CP-element group 311: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_635_loopback_trigger
      -- 
    zeropad_CP_182_elements(311) <= zeropad_CP_182_elements(110);
    -- CP-element group 312:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: successors 
    -- CP-element group 312:  members (2) 
      -- CP-element group 312: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_635_loopback_sample_req
      -- CP-element group 312: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_635_loopback_sample_req_ps
      -- 
    phi_stmt_635_loopback_sample_req_1480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_635_loopback_sample_req_1480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(312), ack => phi_stmt_635_req_0); -- 
    -- Element group zeropad_CP_182_elements(312) is bound as output of CP function.
    -- CP-element group 313:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	111 
    -- CP-element group 313: successors 
    -- CP-element group 313:  members (1) 
      -- CP-element group 313: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_635_entry_trigger
      -- 
    zeropad_CP_182_elements(313) <= zeropad_CP_182_elements(111);
    -- CP-element group 314:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: successors 
    -- CP-element group 314:  members (2) 
      -- CP-element group 314: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_635_entry_sample_req
      -- CP-element group 314: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_635_entry_sample_req_ps
      -- 
    phi_stmt_635_entry_sample_req_1483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_635_entry_sample_req_1483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(314), ack => phi_stmt_635_req_1); -- 
    -- Element group zeropad_CP_182_elements(314) is bound as output of CP function.
    -- CP-element group 315:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: successors 
    -- CP-element group 315:  members (2) 
      -- CP-element group 315: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_635_phi_mux_ack
      -- CP-element group 315: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_635_phi_mux_ack_ps
      -- 
    phi_stmt_635_phi_mux_ack_1486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_635_ack_0, ack => zeropad_CP_182_elements(315)); -- 
    -- CP-element group 316:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	318 
    -- CP-element group 316:  members (1) 
      -- CP-element group 316: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_638_sample_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(316) is bound as output of CP function.
    -- CP-element group 317:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	319 
    -- CP-element group 317:  members (1) 
      -- CP-element group 317: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_638_update_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(317) is bound as output of CP function.
    -- CP-element group 318:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	316 
    -- CP-element group 318: marked-predecessors 
    -- CP-element group 318: 	320 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	320 
    -- CP-element group 318:  members (3) 
      -- CP-element group 318: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_638_sample_start_
      -- CP-element group 318: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_638_Sample/$entry
      -- CP-element group 318: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_638_Sample/rr
      -- 
    rr_1499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(318), ack => type_cast_638_inst_req_0); -- 
    zeropad_cp_element_group_318: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_318"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(316) & zeropad_CP_182_elements(320);
      gj_zeropad_cp_element_group_318 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(318), clk => clk, reset => reset); --
    end block;
    -- CP-element group 319:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	317 
    -- CP-element group 319: marked-predecessors 
    -- CP-element group 319: 	321 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	321 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_638_update_start_
      -- CP-element group 319: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_638_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_638_Update/cr
      -- 
    cr_1504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(319), ack => type_cast_638_inst_req_1); -- 
    zeropad_cp_element_group_319: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_319"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(317) & zeropad_CP_182_elements(321);
      gj_zeropad_cp_element_group_319 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(319), clk => clk, reset => reset); --
    end block;
    -- CP-element group 320:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	318 
    -- CP-element group 320: successors 
    -- CP-element group 320: marked-successors 
    -- CP-element group 320: 	318 
    -- CP-element group 320:  members (4) 
      -- CP-element group 320: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_638_sample_completed__ps
      -- CP-element group 320: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_638_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_638_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_638_Sample/ra
      -- 
    ra_1500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_638_inst_ack_0, ack => zeropad_CP_182_elements(320)); -- 
    -- CP-element group 321:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	319 
    -- CP-element group 321: successors 
    -- CP-element group 321: marked-successors 
    -- CP-element group 321: 	319 
    -- CP-element group 321:  members (4) 
      -- CP-element group 321: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_638_update_completed__ps
      -- CP-element group 321: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_638_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_638_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_638_Update/ca
      -- 
    ca_1505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_638_inst_ack_1, ack => zeropad_CP_182_elements(321)); -- 
    -- CP-element group 322:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: successors 
    -- CP-element group 322:  members (4) 
      -- CP-element group 322: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_valuex_x1_at_entry_639_sample_start__ps
      -- CP-element group 322: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_valuex_x1_at_entry_639_sample_completed__ps
      -- CP-element group 322: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_valuex_x1_at_entry_639_sample_start_
      -- CP-element group 322: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_valuex_x1_at_entry_639_sample_completed_
      -- 
    -- Element group zeropad_CP_182_elements(322) is bound as output of CP function.
    -- CP-element group 323:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	325 
    -- CP-element group 323:  members (2) 
      -- CP-element group 323: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_valuex_x1_at_entry_639_update_start__ps
      -- CP-element group 323: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_valuex_x1_at_entry_639_update_start_
      -- 
    -- Element group zeropad_CP_182_elements(323) is bound as output of CP function.
    -- CP-element group 324:  join  transition  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	325 
    -- CP-element group 324: successors 
    -- CP-element group 324:  members (1) 
      -- CP-element group 324: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_valuex_x1_at_entry_639_update_completed__ps
      -- 
    zeropad_CP_182_elements(324) <= zeropad_CP_182_elements(325);
    -- CP-element group 325:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	323 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	324 
    -- CP-element group 325:  members (1) 
      -- CP-element group 325: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_valuex_x1_at_entry_639_update_completed_
      -- 
    -- Element group zeropad_CP_182_elements(325) is a control-delay.
    cp_element_325_delay: control_delay_element  generic map(name => " 325_delay", delay_value => 1)  port map(req => zeropad_CP_182_elements(323), ack => zeropad_CP_182_elements(325), clk => clk, reset =>reset);
    -- CP-element group 326:  join  transition  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	112 
    -- CP-element group 326: marked-predecessors 
    -- CP-element group 326: 	115 
    -- CP-element group 326: 	401 
    -- CP-element group 326: 	405 
    -- CP-element group 326: 	409 
    -- CP-element group 326: 	521 
    -- CP-element group 326: 	525 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	114 
    -- CP-element group 326:  members (1) 
      -- CP-element group 326: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_640_sample_start_
      -- 
    zeropad_cp_element_group_326: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_326"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(115) & zeropad_CP_182_elements(401) & zeropad_CP_182_elements(405) & zeropad_CP_182_elements(409) & zeropad_CP_182_elements(521) & zeropad_CP_182_elements(525);
      gj_zeropad_cp_element_group_326 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(326), clk => clk, reset => reset); --
    end block;
    -- CP-element group 327:  join  transition  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	112 
    -- CP-element group 327: marked-predecessors 
    -- CP-element group 327: 	331 
    -- CP-element group 327: 	373 
    -- CP-element group 327: 	408 
    -- CP-element group 327: 	524 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	116 
    -- CP-element group 327:  members (1) 
      -- CP-element group 327: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_640_update_start_
      -- 
    zeropad_cp_element_group_327: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_327"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(331) & zeropad_CP_182_elements(373) & zeropad_CP_182_elements(408) & zeropad_CP_182_elements(524);
      gj_zeropad_cp_element_group_327 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(327), clk => clk, reset => reset); --
    end block;
    -- CP-element group 328:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	114 
    -- CP-element group 328: successors 
    -- CP-element group 328:  members (1) 
      -- CP-element group 328: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_640_sample_start__ps
      -- 
    zeropad_CP_182_elements(328) <= zeropad_CP_182_elements(114);
    -- CP-element group 329:  join  transition  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	115 
    -- CP-element group 329:  members (1) 
      -- CP-element group 329: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_640_sample_completed__ps
      -- 
    -- Element group zeropad_CP_182_elements(329) is bound as output of CP function.
    -- CP-element group 330:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	116 
    -- CP-element group 330: successors 
    -- CP-element group 330:  members (1) 
      -- CP-element group 330: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_640_update_start__ps
      -- 
    zeropad_CP_182_elements(330) <= zeropad_CP_182_elements(116);
    -- CP-element group 331:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	117 
    -- CP-element group 331: 	371 
    -- CP-element group 331: 	406 
    -- CP-element group 331: 	522 
    -- CP-element group 331: marked-successors 
    -- CP-element group 331: 	327 
    -- CP-element group 331:  members (2) 
      -- CP-element group 331: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_640_update_completed_
      -- CP-element group 331: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_640_update_completed__ps
      -- 
    -- Element group zeropad_CP_182_elements(331) is bound as output of CP function.
    -- CP-element group 332:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	110 
    -- CP-element group 332: successors 
    -- CP-element group 332:  members (1) 
      -- CP-element group 332: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_640_loopback_trigger
      -- 
    zeropad_CP_182_elements(332) <= zeropad_CP_182_elements(110);
    -- CP-element group 333:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: successors 
    -- CP-element group 333:  members (2) 
      -- CP-element group 333: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_640_loopback_sample_req
      -- CP-element group 333: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_640_loopback_sample_req_ps
      -- 
    phi_stmt_640_loopback_sample_req_1524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_640_loopback_sample_req_1524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(333), ack => phi_stmt_640_req_0); -- 
    -- Element group zeropad_CP_182_elements(333) is bound as output of CP function.
    -- CP-element group 334:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	111 
    -- CP-element group 334: successors 
    -- CP-element group 334:  members (1) 
      -- CP-element group 334: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_640_entry_trigger
      -- 
    zeropad_CP_182_elements(334) <= zeropad_CP_182_elements(111);
    -- CP-element group 335:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: successors 
    -- CP-element group 335:  members (2) 
      -- CP-element group 335: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_640_entry_sample_req
      -- CP-element group 335: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_640_entry_sample_req_ps
      -- 
    phi_stmt_640_entry_sample_req_1527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_640_entry_sample_req_1527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(335), ack => phi_stmt_640_req_1); -- 
    -- Element group zeropad_CP_182_elements(335) is bound as output of CP function.
    -- CP-element group 336:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: successors 
    -- CP-element group 336:  members (2) 
      -- CP-element group 336: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_640_phi_mux_ack
      -- CP-element group 336: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/phi_stmt_640_phi_mux_ack_ps
      -- 
    phi_stmt_640_phi_mux_ack_1530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_640_ack_0, ack => zeropad_CP_182_elements(336)); -- 
    -- CP-element group 337:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	339 
    -- CP-element group 337:  members (1) 
      -- CP-element group 337: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_643_sample_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(337) is bound as output of CP function.
    -- CP-element group 338:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	340 
    -- CP-element group 338:  members (1) 
      -- CP-element group 338: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_643_update_start__ps
      -- 
    -- Element group zeropad_CP_182_elements(338) is bound as output of CP function.
    -- CP-element group 339:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	337 
    -- CP-element group 339: marked-predecessors 
    -- CP-element group 339: 	341 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	341 
    -- CP-element group 339:  members (3) 
      -- CP-element group 339: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_643_sample_start_
      -- CP-element group 339: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_643_Sample/$entry
      -- CP-element group 339: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_643_Sample/rr
      -- 
    rr_1543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(339), ack => type_cast_643_inst_req_0); -- 
    zeropad_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(337) & zeropad_CP_182_elements(341);
      gj_zeropad_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: marked-predecessors 
    -- CP-element group 340: 	342 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	342 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_643_update_start_
      -- CP-element group 340: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_643_Update/$entry
      -- CP-element group 340: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_643_Update/cr
      -- 
    cr_1548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(340), ack => type_cast_643_inst_req_1); -- 
    zeropad_cp_element_group_340: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_340"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(338) & zeropad_CP_182_elements(342);
      gj_zeropad_cp_element_group_340 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(340), clk => clk, reset => reset); --
    end block;
    -- CP-element group 341:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	339 
    -- CP-element group 341: successors 
    -- CP-element group 341: marked-successors 
    -- CP-element group 341: 	339 
    -- CP-element group 341:  members (4) 
      -- CP-element group 341: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_643_sample_completed__ps
      -- CP-element group 341: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_643_sample_completed_
      -- CP-element group 341: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_643_Sample/$exit
      -- CP-element group 341: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_643_Sample/ra
      -- 
    ra_1544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_643_inst_ack_0, ack => zeropad_CP_182_elements(341)); -- 
    -- CP-element group 342:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	340 
    -- CP-element group 342: successors 
    -- CP-element group 342: marked-successors 
    -- CP-element group 342: 	340 
    -- CP-element group 342:  members (4) 
      -- CP-element group 342: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_643_update_completed__ps
      -- CP-element group 342: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_643_update_completed_
      -- CP-element group 342: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_643_Update/$exit
      -- CP-element group 342: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_643_Update/ca
      -- 
    ca_1549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_643_inst_ack_1, ack => zeropad_CP_182_elements(342)); -- 
    -- CP-element group 343:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	345 
    -- CP-element group 343:  members (4) 
      -- CP-element group 343: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_wordx_x1_at_entry_644_sample_start__ps
      -- CP-element group 343: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_wordx_x1_at_entry_644_sample_start_
      -- CP-element group 343: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_wordx_x1_at_entry_644_Sample/$entry
      -- CP-element group 343: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_wordx_x1_at_entry_644_Sample/req
      -- 
    req_1561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(343), ack => input_wordx_x1_at_entry_583_644_buf_req_0); -- 
    -- Element group zeropad_CP_182_elements(343) is bound as output of CP function.
    -- CP-element group 344:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	346 
    -- CP-element group 344:  members (4) 
      -- CP-element group 344: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_wordx_x1_at_entry_644_update_start__ps
      -- CP-element group 344: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_wordx_x1_at_entry_644_update_start_
      -- CP-element group 344: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_wordx_x1_at_entry_644_Update/$entry
      -- CP-element group 344: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_wordx_x1_at_entry_644_Update/req
      -- 
    req_1566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(344), ack => input_wordx_x1_at_entry_583_644_buf_req_1); -- 
    -- Element group zeropad_CP_182_elements(344) is bound as output of CP function.
    -- CP-element group 345:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	343 
    -- CP-element group 345: successors 
    -- CP-element group 345:  members (4) 
      -- CP-element group 345: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_wordx_x1_at_entry_644_sample_completed__ps
      -- CP-element group 345: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_wordx_x1_at_entry_644_sample_completed_
      -- CP-element group 345: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_wordx_x1_at_entry_644_Sample/$exit
      -- CP-element group 345: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_wordx_x1_at_entry_644_Sample/ack
      -- 
    ack_1562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => input_wordx_x1_at_entry_583_644_buf_ack_0, ack => zeropad_CP_182_elements(345)); -- 
    -- CP-element group 346:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	344 
    -- CP-element group 346: successors 
    -- CP-element group 346:  members (4) 
      -- CP-element group 346: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_wordx_x1_at_entry_644_update_completed__ps
      -- CP-element group 346: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_wordx_x1_at_entry_644_update_completed_
      -- CP-element group 346: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_wordx_x1_at_entry_644_Update/$exit
      -- CP-element group 346: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/R_input_wordx_x1_at_entry_644_Update/ack
      -- 
    ack_1567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => input_wordx_x1_at_entry_583_644_buf_ack_1, ack => zeropad_CP_182_elements(346)); -- 
    -- CP-element group 347:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	142 
    -- CP-element group 347: 	163 
    -- CP-element group 347: 	226 
    -- CP-element group 347: marked-predecessors 
    -- CP-element group 347: 	349 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	349 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_684_sample_start_
      -- CP-element group 347: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_684_Sample/$entry
      -- CP-element group 347: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_684_Sample/rr
      -- 
    rr_1576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(347), ack => type_cast_684_inst_req_0); -- 
    zeropad_cp_element_group_347: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_347"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(226) & zeropad_CP_182_elements(349);
      gj_zeropad_cp_element_group_347 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(347), clk => clk, reset => reset); --
    end block;
    -- CP-element group 348:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: marked-predecessors 
    -- CP-element group 348: 	350 
    -- CP-element group 348: 	365 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	350 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_684_update_start_
      -- CP-element group 348: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_684_Update/$entry
      -- CP-element group 348: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_684_Update/cr
      -- 
    cr_1581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(348), ack => type_cast_684_inst_req_1); -- 
    zeropad_cp_element_group_348: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_348"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(350) & zeropad_CP_182_elements(365);
      gj_zeropad_cp_element_group_348 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(348), clk => clk, reset => reset); --
    end block;
    -- CP-element group 349:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	347 
    -- CP-element group 349: successors 
    -- CP-element group 349: marked-successors 
    -- CP-element group 349: 	138 
    -- CP-element group 349: 	159 
    -- CP-element group 349: 	222 
    -- CP-element group 349: 	347 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_684_sample_completed_
      -- CP-element group 349: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_684_Sample/$exit
      -- CP-element group 349: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_684_Sample/ra
      -- 
    ra_1577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_684_inst_ack_0, ack => zeropad_CP_182_elements(349)); -- 
    -- CP-element group 350:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	348 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	363 
    -- CP-element group 350: marked-successors 
    -- CP-element group 350: 	348 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_684_update_completed_
      -- CP-element group 350: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_684_Update/$exit
      -- CP-element group 350: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_684_Update/ca
      -- 
    ca_1582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_684_inst_ack_1, ack => zeropad_CP_182_elements(350)); -- 
    -- CP-element group 351:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	142 
    -- CP-element group 351: 	163 
    -- CP-element group 351: marked-predecessors 
    -- CP-element group 351: 	353 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	353 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_688_sample_start_
      -- CP-element group 351: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_688_Sample/$entry
      -- CP-element group 351: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_688_Sample/req
      -- 
    req_1590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(351), ack => W_ifx_xend_exec_guard_686_delayed_1_0_686_inst_req_0); -- 
    zeropad_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(353);
      gj_zeropad_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: marked-predecessors 
    -- CP-element group 352: 	354 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	354 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_688_update_start_
      -- CP-element group 352: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_688_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_688_Update/req
      -- 
    req_1595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(352), ack => W_ifx_xend_exec_guard_686_delayed_1_0_686_inst_req_1); -- 
    zeropad_cp_element_group_352: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_352"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_CP_182_elements(354);
      gj_zeropad_cp_element_group_352 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(352), clk => clk, reset => reset); --
    end block;
    -- CP-element group 353:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	351 
    -- CP-element group 353: successors 
    -- CP-element group 353: marked-successors 
    -- CP-element group 353: 	138 
    -- CP-element group 353: 	159 
    -- CP-element group 353: 	351 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_688_sample_completed_
      -- CP-element group 353: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_688_Sample/$exit
      -- CP-element group 353: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_688_Sample/ack
      -- 
    ack_1591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_686_delayed_1_0_686_inst_ack_0, ack => zeropad_CP_182_elements(353)); -- 
    -- CP-element group 354:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	352 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	611 
    -- CP-element group 354: marked-successors 
    -- CP-element group 354: 	352 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_688_update_completed_
      -- CP-element group 354: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_688_Update/$exit
      -- CP-element group 354: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_688_Update/ack
      -- 
    ack_1596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_686_delayed_1_0_686_inst_ack_1, ack => zeropad_CP_182_elements(354)); -- 
    -- CP-element group 355:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	142 
    -- CP-element group 355: 	163 
    -- CP-element group 355: marked-predecessors 
    -- CP-element group 355: 	357 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	357 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_698_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_698_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_698_Sample/req
      -- 
    req_1604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(355), ack => W_ifx_xend_exec_guard_693_delayed_1_0_696_inst_req_0); -- 
    zeropad_cp_element_group_355: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_355"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(357);
      gj_zeropad_cp_element_group_355 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(355), clk => clk, reset => reset); --
    end block;
    -- CP-element group 356:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: marked-predecessors 
    -- CP-element group 356: 	358 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	358 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_698_update_start_
      -- CP-element group 356: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_698_Update/$entry
      -- CP-element group 356: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_698_Update/req
      -- 
    req_1609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(356), ack => W_ifx_xend_exec_guard_693_delayed_1_0_696_inst_req_1); -- 
    zeropad_cp_element_group_356: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_356"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_CP_182_elements(358);
      gj_zeropad_cp_element_group_356 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(356), clk => clk, reset => reset); --
    end block;
    -- CP-element group 357:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	355 
    -- CP-element group 357: successors 
    -- CP-element group 357: marked-successors 
    -- CP-element group 357: 	138 
    -- CP-element group 357: 	159 
    -- CP-element group 357: 	355 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_698_sample_completed_
      -- CP-element group 357: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_698_Sample/$exit
      -- CP-element group 357: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_698_Sample/ack
      -- 
    ack_1605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_693_delayed_1_0_696_inst_ack_0, ack => zeropad_CP_182_elements(357)); -- 
    -- CP-element group 358:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	356 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	611 
    -- CP-element group 358: marked-successors 
    -- CP-element group 358: 	356 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_698_update_completed_
      -- CP-element group 358: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_698_Update/$exit
      -- CP-element group 358: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_698_Update/ack
      -- 
    ack_1610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_693_delayed_1_0_696_inst_ack_1, ack => zeropad_CP_182_elements(358)); -- 
    -- CP-element group 359:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	142 
    -- CP-element group 359: 	163 
    -- CP-element group 359: marked-predecessors 
    -- CP-element group 359: 	361 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	361 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_708_sample_start_
      -- CP-element group 359: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_708_Sample/$entry
      -- CP-element group 359: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_708_Sample/req
      -- 
    req_1618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(359), ack => W_ifx_xend_exec_guard_700_delayed_1_0_706_inst_req_0); -- 
    zeropad_cp_element_group_359: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_359"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(361);
      gj_zeropad_cp_element_group_359 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(359), clk => clk, reset => reset); --
    end block;
    -- CP-element group 360:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: marked-predecessors 
    -- CP-element group 360: 	362 
    -- CP-element group 360: 	365 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	362 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_708_update_start_
      -- CP-element group 360: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_708_Update/$entry
      -- CP-element group 360: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_708_Update/req
      -- 
    req_1623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(360), ack => W_ifx_xend_exec_guard_700_delayed_1_0_706_inst_req_1); -- 
    zeropad_cp_element_group_360: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_360"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(362) & zeropad_CP_182_elements(365);
      gj_zeropad_cp_element_group_360 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(360), clk => clk, reset => reset); --
    end block;
    -- CP-element group 361:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	359 
    -- CP-element group 361: successors 
    -- CP-element group 361: marked-successors 
    -- CP-element group 361: 	138 
    -- CP-element group 361: 	159 
    -- CP-element group 361: 	359 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_708_sample_completed_
      -- CP-element group 361: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_708_Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_708_Sample/ack
      -- 
    ack_1619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_700_delayed_1_0_706_inst_ack_0, ack => zeropad_CP_182_elements(361)); -- 
    -- CP-element group 362:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	360 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362: marked-successors 
    -- CP-element group 362: 	360 
    -- CP-element group 362:  members (3) 
      -- CP-element group 362: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_708_update_completed_
      -- CP-element group 362: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_708_Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_708_Update/ack
      -- 
    ack_1624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_700_delayed_1_0_706_inst_ack_1, ack => zeropad_CP_182_elements(362)); -- 
    -- CP-element group 363:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	350 
    -- CP-element group 363: 	362 
    -- CP-element group 363: marked-predecessors 
    -- CP-element group 363: 	365 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	365 
    -- CP-element group 363:  members (3) 
      -- CP-element group 363: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_712_sample_start_
      -- CP-element group 363: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_712_Sample/$entry
      -- CP-element group 363: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_712_Sample/rr
      -- 
    rr_1632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(363), ack => type_cast_712_inst_req_0); -- 
    zeropad_cp_element_group_363: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_363"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(350) & zeropad_CP_182_elements(362) & zeropad_CP_182_elements(365);
      gj_zeropad_cp_element_group_363 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(363), clk => clk, reset => reset); --
    end block;
    -- CP-element group 364:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	115 
    -- CP-element group 364: marked-predecessors 
    -- CP-element group 364: 	366 
    -- CP-element group 364: 	571 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	366 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_712_update_start_
      -- CP-element group 364: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_712_Update/$entry
      -- CP-element group 364: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_712_Update/cr
      -- 
    cr_1637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(364), ack => type_cast_712_inst_req_1); -- 
    zeropad_cp_element_group_364: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_364"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(366) & zeropad_CP_182_elements(571);
      gj_zeropad_cp_element_group_364 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(364), clk => clk, reset => reset); --
    end block;
    -- CP-element group 365:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	363 
    -- CP-element group 365: successors 
    -- CP-element group 365: marked-successors 
    -- CP-element group 365: 	348 
    -- CP-element group 365: 	360 
    -- CP-element group 365: 	363 
    -- CP-element group 365:  members (3) 
      -- CP-element group 365: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_712_sample_completed_
      -- CP-element group 365: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_712_Sample/$exit
      -- CP-element group 365: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_712_Sample/ra
      -- 
    ra_1633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_712_inst_ack_0, ack => zeropad_CP_182_elements(365)); -- 
    -- CP-element group 366:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	364 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	569 
    -- CP-element group 366: marked-successors 
    -- CP-element group 366: 	305 
    -- CP-element group 366: 	364 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_712_update_completed_
      -- CP-element group 366: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_712_Update/$exit
      -- CP-element group 366: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_712_Update/ca
      -- 
    ca_1638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_712_inst_ack_1, ack => zeropad_CP_182_elements(366)); -- 
    -- CP-element group 367:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	142 
    -- CP-element group 367: 	163 
    -- CP-element group 367: marked-predecessors 
    -- CP-element group 367: 	369 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	369 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_716_sample_start_
      -- CP-element group 367: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_716_Sample/$entry
      -- CP-element group 367: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_716_Sample/req
      -- 
    req_1646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(367), ack => W_ifx_xend_exec_guard_705_delayed_2_0_714_inst_req_0); -- 
    zeropad_cp_element_group_367: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_367"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(369);
      gj_zeropad_cp_element_group_367 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(367), clk => clk, reset => reset); --
    end block;
    -- CP-element group 368:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: marked-predecessors 
    -- CP-element group 368: 	370 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	370 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_716_update_start_
      -- CP-element group 368: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_716_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_716_Update/req
      -- 
    req_1651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(368), ack => W_ifx_xend_exec_guard_705_delayed_2_0_714_inst_req_1); -- 
    zeropad_cp_element_group_368: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_368"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_CP_182_elements(370);
      gj_zeropad_cp_element_group_368 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(368), clk => clk, reset => reset); --
    end block;
    -- CP-element group 369:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	367 
    -- CP-element group 369: successors 
    -- CP-element group 369: marked-successors 
    -- CP-element group 369: 	138 
    -- CP-element group 369: 	159 
    -- CP-element group 369: 	367 
    -- CP-element group 369:  members (3) 
      -- CP-element group 369: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_716_sample_completed_
      -- CP-element group 369: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_716_Sample/$exit
      -- CP-element group 369: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_716_Sample/ack
      -- 
    ack_1647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_705_delayed_2_0_714_inst_ack_0, ack => zeropad_CP_182_elements(369)); -- 
    -- CP-element group 370:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	368 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	611 
    -- CP-element group 370: marked-successors 
    -- CP-element group 370: 	368 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_716_update_completed_
      -- CP-element group 370: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_716_Update/$exit
      -- CP-element group 370: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_716_Update/ack
      -- 
    ack_1652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_705_delayed_2_0_714_inst_ack_1, ack => zeropad_CP_182_elements(370)); -- 
    -- CP-element group 371:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	331 
    -- CP-element group 371: marked-predecessors 
    -- CP-element group 371: 	373 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	373 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_719_sample_start_
      -- CP-element group 371: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_719_Sample/$entry
      -- CP-element group 371: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_719_Sample/req
      -- 
    req_1660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(371), ack => W_input_wordx_x1_707_delayed_2_0_717_inst_req_0); -- 
    zeropad_cp_element_group_371: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_371"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(331) & zeropad_CP_182_elements(373);
      gj_zeropad_cp_element_group_371 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(371), clk => clk, reset => reset); --
    end block;
    -- CP-element group 372:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	115 
    -- CP-element group 372: marked-predecessors 
    -- CP-element group 372: 	374 
    -- CP-element group 372: 	571 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	374 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_719_update_start_
      -- CP-element group 372: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_719_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_719_Update/req
      -- 
    req_1665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(372), ack => W_input_wordx_x1_707_delayed_2_0_717_inst_req_1); -- 
    zeropad_cp_element_group_372: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_372"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(374) & zeropad_CP_182_elements(571);
      gj_zeropad_cp_element_group_372 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(372), clk => clk, reset => reset); --
    end block;
    -- CP-element group 373:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	371 
    -- CP-element group 373: successors 
    -- CP-element group 373: marked-successors 
    -- CP-element group 373: 	327 
    -- CP-element group 373: 	371 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_719_sample_completed_
      -- CP-element group 373: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_719_Sample/$exit
      -- CP-element group 373: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_719_Sample/ack
      -- 
    ack_1661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_wordx_x1_707_delayed_2_0_717_inst_ack_0, ack => zeropad_CP_182_elements(373)); -- 
    -- CP-element group 374:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	372 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	569 
    -- CP-element group 374: marked-successors 
    -- CP-element group 374: 	305 
    -- CP-element group 374: 	372 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_719_update_completed_
      -- CP-element group 374: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_719_Update/$exit
      -- CP-element group 374: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_719_Update/ack
      -- 
    ack_1666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_input_wordx_x1_707_delayed_2_0_717_inst_ack_1, ack => zeropad_CP_182_elements(374)); -- 
    -- CP-element group 375:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	142 
    -- CP-element group 375: 	163 
    -- CP-element group 375: marked-predecessors 
    -- CP-element group 375: 	377 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	377 
    -- CP-element group 375:  members (3) 
      -- CP-element group 375: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_735_sample_start_
      -- CP-element group 375: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_735_Sample/$entry
      -- CP-element group 375: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_735_Sample/req
      -- 
    req_1674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(375), ack => W_ifx_xend_exec_guard_718_delayed_2_0_733_inst_req_0); -- 
    zeropad_cp_element_group_375: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_375"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(377);
      gj_zeropad_cp_element_group_375 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(375), clk => clk, reset => reset); --
    end block;
    -- CP-element group 376:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: marked-predecessors 
    -- CP-element group 376: 	378 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	378 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_735_update_start_
      -- CP-element group 376: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_735_Update/$entry
      -- CP-element group 376: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_735_Update/req
      -- 
    req_1679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(376), ack => W_ifx_xend_exec_guard_718_delayed_2_0_733_inst_req_1); -- 
    zeropad_cp_element_group_376: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_376"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_CP_182_elements(378);
      gj_zeropad_cp_element_group_376 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(376), clk => clk, reset => reset); --
    end block;
    -- CP-element group 377:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	375 
    -- CP-element group 377: successors 
    -- CP-element group 377: marked-successors 
    -- CP-element group 377: 	138 
    -- CP-element group 377: 	159 
    -- CP-element group 377: 	375 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_735_sample_completed_
      -- CP-element group 377: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_735_Sample/$exit
      -- CP-element group 377: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_735_Sample/ack
      -- 
    ack_1675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_718_delayed_2_0_733_inst_ack_0, ack => zeropad_CP_182_elements(377)); -- 
    -- CP-element group 378:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	376 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	611 
    -- CP-element group 378: marked-successors 
    -- CP-element group 378: 	376 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_735_update_completed_
      -- CP-element group 378: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_735_Update/$exit
      -- CP-element group 378: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_735_Update/ack
      -- 
    ack_1680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_718_delayed_2_0_733_inst_ack_1, ack => zeropad_CP_182_elements(378)); -- 
    -- CP-element group 379:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	142 
    -- CP-element group 379: 	163 
    -- CP-element group 379: marked-predecessors 
    -- CP-element group 379: 	381 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	381 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_745_sample_start_
      -- CP-element group 379: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_745_Sample/$entry
      -- CP-element group 379: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_745_Sample/req
      -- 
    req_1688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(379), ack => W_ifx_xend_exec_guard_725_delayed_2_0_743_inst_req_0); -- 
    zeropad_cp_element_group_379: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_379"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(381);
      gj_zeropad_cp_element_group_379 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(379), clk => clk, reset => reset); --
    end block;
    -- CP-element group 380:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: marked-predecessors 
    -- CP-element group 380: 	382 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	382 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_745_update_start_
      -- CP-element group 380: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_745_Update/$entry
      -- CP-element group 380: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_745_Update/req
      -- 
    req_1693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(380), ack => W_ifx_xend_exec_guard_725_delayed_2_0_743_inst_req_1); -- 
    zeropad_cp_element_group_380: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_380"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_CP_182_elements(382);
      gj_zeropad_cp_element_group_380 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(380), clk => clk, reset => reset); --
    end block;
    -- CP-element group 381:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	379 
    -- CP-element group 381: successors 
    -- CP-element group 381: marked-successors 
    -- CP-element group 381: 	138 
    -- CP-element group 381: 	159 
    -- CP-element group 381: 	379 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_745_sample_completed_
      -- CP-element group 381: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_745_Sample/$exit
      -- CP-element group 381: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_745_Sample/ack
      -- 
    ack_1689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_725_delayed_2_0_743_inst_ack_0, ack => zeropad_CP_182_elements(381)); -- 
    -- CP-element group 382:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	380 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	611 
    -- CP-element group 382: marked-successors 
    -- CP-element group 382: 	380 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_745_update_completed_
      -- CP-element group 382: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_745_Update/$exit
      -- CP-element group 382: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_745_Update/ack
      -- 
    ack_1694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend_exec_guard_725_delayed_2_0_743_inst_ack_1, ack => zeropad_CP_182_elements(382)); -- 
    -- CP-element group 383:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	310 
    -- CP-element group 383: marked-predecessors 
    -- CP-element group 383: 	385 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	385 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_748_sample_start_
      -- CP-element group 383: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_748_Sample/$entry
      -- CP-element group 383: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_748_Sample/req
      -- 
    req_1702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(383), ack => W_shl169_728_delayed_2_0_746_inst_req_0); -- 
    zeropad_cp_element_group_383: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_383"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(310) & zeropad_CP_182_elements(385);
      gj_zeropad_cp_element_group_383 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(383), clk => clk, reset => reset); --
    end block;
    -- CP-element group 384:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	115 
    -- CP-element group 384: marked-predecessors 
    -- CP-element group 384: 	386 
    -- CP-element group 384: 	571 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	386 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_748_update_start_
      -- CP-element group 384: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_748_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_748_Update/req
      -- 
    req_1707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(384), ack => W_shl169_728_delayed_2_0_746_inst_req_1); -- 
    zeropad_cp_element_group_384: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_384"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(386) & zeropad_CP_182_elements(571);
      gj_zeropad_cp_element_group_384 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(384), clk => clk, reset => reset); --
    end block;
    -- CP-element group 385:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	383 
    -- CP-element group 385: successors 
    -- CP-element group 385: marked-successors 
    -- CP-element group 385: 	306 
    -- CP-element group 385: 	383 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_748_sample_completed_
      -- CP-element group 385: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_748_Sample/$exit
      -- CP-element group 385: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_748_Sample/ack
      -- 
    ack_1703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 385_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_shl169_728_delayed_2_0_746_inst_ack_0, ack => zeropad_CP_182_elements(385)); -- 
    -- CP-element group 386:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	384 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	569 
    -- CP-element group 386: marked-successors 
    -- CP-element group 386: 	305 
    -- CP-element group 386: 	384 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_748_update_completed_
      -- CP-element group 386: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_748_Update/$exit
      -- CP-element group 386: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_748_Update/ack
      -- 
    ack_1708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_shl169_728_delayed_2_0_746_inst_ack_1, ack => zeropad_CP_182_elements(386)); -- 
    -- CP-element group 387:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	391 
    -- CP-element group 387: marked-predecessors 
    -- CP-element group 387: 	392 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	392 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_790_request/req
      -- CP-element group 387: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_790_request/$entry
      -- CP-element group 387: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_790_sample_start_
      -- 
    req_1748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(387), ack => addr_of_790_final_reg_req_0); -- 
    zeropad_cp_element_group_387: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_387"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(391) & zeropad_CP_182_elements(392);
      gj_zeropad_cp_element_group_387 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(387), clk => clk, reset => reset); --
    end block;
    -- CP-element group 388:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	112 
    -- CP-element group 388: marked-predecessors 
    -- CP-element group 388: 	393 
    -- CP-element group 388: 	400 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	393 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_790_complete/req
      -- CP-element group 388: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_790_complete/$entry
      -- CP-element group 388: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_790_update_start_
      -- 
    req_1753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(388), ack => addr_of_790_final_reg_req_1); -- 
    zeropad_cp_element_group_388: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_388"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(393) & zeropad_CP_182_elements(400);
      gj_zeropad_cp_element_group_388 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(388), clk => clk, reset => reset); --
    end block;
    -- CP-element group 389:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	112 
    -- CP-element group 389: marked-predecessors 
    -- CP-element group 389: 	391 
    -- CP-element group 389: 	392 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	391 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_final_index_sum_regn_Update/$entry
      -- CP-element group 389: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_final_index_sum_regn_update_start
      -- CP-element group 389: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_final_index_sum_regn_Update/req
      -- 
    req_1738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(389), ack => array_obj_ref_789_index_offset_req_1); -- 
    zeropad_cp_element_group_389: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_389"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(391) & zeropad_CP_182_elements(392);
      gj_zeropad_cp_element_group_389 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(389), clk => clk, reset => reset); --
    end block;
    -- CP-element group 390:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	121 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	611 
    -- CP-element group 390: marked-successors 
    -- CP-element group 390: 	119 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_final_index_sum_regn_Sample/ack
      -- CP-element group 390: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_final_index_sum_regn_Sample/$exit
      -- CP-element group 390: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_final_index_sum_regn_sample_complete
      -- 
    ack_1734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_789_index_offset_ack_0, ack => zeropad_CP_182_elements(390)); -- 
    -- CP-element group 391:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	389 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	387 
    -- CP-element group 391: marked-successors 
    -- CP-element group 391: 	389 
    -- CP-element group 391:  members (8) 
      -- CP-element group 391: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_final_index_sum_regn_Update/ack
      -- CP-element group 391: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_base_plus_offset/$entry
      -- CP-element group 391: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_base_plus_offset/$exit
      -- CP-element group 391: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_base_plus_offset/sum_rename_ack
      -- CP-element group 391: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_final_index_sum_regn_Update/$exit
      -- CP-element group 391: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_base_plus_offset/sum_rename_req
      -- CP-element group 391: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_root_address_calculated
      -- CP-element group 391: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_789_offset_calculated
      -- 
    ack_1739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_789_index_offset_ack_1, ack => zeropad_CP_182_elements(391)); -- 
    -- CP-element group 392:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	387 
    -- CP-element group 392: successors 
    -- CP-element group 392: marked-successors 
    -- CP-element group 392: 	387 
    -- CP-element group 392: 	389 
    -- CP-element group 392:  members (3) 
      -- CP-element group 392: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_790_request/$exit
      -- CP-element group 392: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_790_request/ack
      -- CP-element group 392: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_790_sample_completed_
      -- 
    ack_1749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_790_final_reg_ack_0, ack => zeropad_CP_182_elements(392)); -- 
    -- CP-element group 393:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	388 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	398 
    -- CP-element group 393: marked-successors 
    -- CP-element group 393: 	388 
    -- CP-element group 393:  members (19) 
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_root_address_calculated
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_base_addr_resize/base_resize_req
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_word_address_calculated
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_base_addr_resize/$exit
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_790_complete/$exit
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_base_plus_offset/sum_rename_req
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_base_plus_offset/sum_rename_ack
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_base_address_resized
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_base_plus_offset/$entry
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_word_addrgen/$entry
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_base_addr_resize/$entry
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_word_addrgen/root_register_req
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_word_addrgen/$exit
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_base_addr_resize/base_resize_ack
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_base_plus_offset/$exit
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_base_address_calculated
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_790_complete/ack
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_word_addrgen/root_register_ack
      -- CP-element group 393: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_790_update_completed_
      -- 
    ack_1754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_790_final_reg_ack_1, ack => zeropad_CP_182_elements(393)); -- 
    -- CP-element group 394:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	142 
    -- CP-element group 394: 	163 
    -- CP-element group 394: 	226 
    -- CP-element group 394: marked-predecessors 
    -- CP-element group 394: 	396 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	396 
    -- CP-element group 394:  members (3) 
      -- CP-element group 394: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_794_sample_start_
      -- CP-element group 394: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_794_Sample/$entry
      -- CP-element group 394: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_794_Sample/req
      -- 
    req_1762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(394), ack => W_ifx_xthen180_exec_guard_768_delayed_6_0_792_inst_req_0); -- 
    zeropad_cp_element_group_394: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_394"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(226) & zeropad_CP_182_elements(396);
      gj_zeropad_cp_element_group_394 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(394), clk => clk, reset => reset); --
    end block;
    -- CP-element group 395:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: marked-predecessors 
    -- CP-element group 395: 	397 
    -- CP-element group 395: 	400 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	397 
    -- CP-element group 395:  members (3) 
      -- CP-element group 395: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_794_update_start_
      -- CP-element group 395: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_794_Update/$entry
      -- CP-element group 395: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_794_Update/req
      -- 
    req_1767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(395), ack => W_ifx_xthen180_exec_guard_768_delayed_6_0_792_inst_req_1); -- 
    zeropad_cp_element_group_395: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_395"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(397) & zeropad_CP_182_elements(400);
      gj_zeropad_cp_element_group_395 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(395), clk => clk, reset => reset); --
    end block;
    -- CP-element group 396:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	394 
    -- CP-element group 396: successors 
    -- CP-element group 396: marked-successors 
    -- CP-element group 396: 	138 
    -- CP-element group 396: 	159 
    -- CP-element group 396: 	222 
    -- CP-element group 396: 	394 
    -- CP-element group 396:  members (3) 
      -- CP-element group 396: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_794_sample_completed_
      -- CP-element group 396: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_794_Sample/$exit
      -- CP-element group 396: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_794_Sample/ack
      -- 
    ack_1763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen180_exec_guard_768_delayed_6_0_792_inst_ack_0, ack => zeropad_CP_182_elements(396)); -- 
    -- CP-element group 397:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	395 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	398 
    -- CP-element group 397: marked-successors 
    -- CP-element group 397: 	395 
    -- CP-element group 397:  members (3) 
      -- CP-element group 397: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_794_update_completed_
      -- CP-element group 397: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_794_Update/$exit
      -- CP-element group 397: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_794_Update/ack
      -- 
    ack_1768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen180_exec_guard_768_delayed_6_0_792_inst_ack_1, ack => zeropad_CP_182_elements(397)); -- 
    -- CP-element group 398:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	393 
    -- CP-element group 398: 	397 
    -- CP-element group 398: marked-predecessors 
    -- CP-element group 398: 	400 
    -- CP-element group 398: 	571 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	400 
    -- CP-element group 398:  members (5) 
      -- CP-element group 398: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_sample_start_
      -- CP-element group 398: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Sample/$entry
      -- CP-element group 398: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Sample/word_access_start/$entry
      -- CP-element group 398: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Sample/word_access_start/word_0/$entry
      -- CP-element group 398: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Sample/word_access_start/word_0/rr
      -- 
    rr_1801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(398), ack => ptr_deref_798_load_0_req_0); -- 
    zeropad_cp_element_group_398: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_398"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(393) & zeropad_CP_182_elements(397) & zeropad_CP_182_elements(400) & zeropad_CP_182_elements(571);
      gj_zeropad_cp_element_group_398 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(398), clk => clk, reset => reset); --
    end block;
    -- CP-element group 399:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	115 
    -- CP-element group 399: marked-predecessors 
    -- CP-element group 399: 	401 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	401 
    -- CP-element group 399:  members (5) 
      -- CP-element group 399: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_update_start_
      -- CP-element group 399: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Update/word_access_complete/word_0/cr
      -- CP-element group 399: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Update/word_access_complete/$entry
      -- CP-element group 399: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Update/word_access_complete/word_0/$entry
      -- 
    cr_1812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(399), ack => ptr_deref_798_load_0_req_1); -- 
    zeropad_cp_element_group_399: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_399"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(401);
      gj_zeropad_cp_element_group_399 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(399), clk => clk, reset => reset); --
    end block;
    -- CP-element group 400:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	398 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	610 
    -- CP-element group 400: marked-successors 
    -- CP-element group 400: 	388 
    -- CP-element group 400: 	395 
    -- CP-element group 400: 	398 
    -- CP-element group 400:  members (5) 
      -- CP-element group 400: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_sample_completed_
      -- CP-element group 400: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Sample/$exit
      -- CP-element group 400: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Sample/word_access_start/$exit
      -- CP-element group 400: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Sample/word_access_start/word_0/$exit
      -- CP-element group 400: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Sample/word_access_start/word_0/ra
      -- 
    ra_1802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_798_load_0_ack_0, ack => zeropad_CP_182_elements(400)); -- 
    -- CP-element group 401:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	399 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	611 
    -- CP-element group 401: marked-successors 
    -- CP-element group 401: 	326 
    -- CP-element group 401: 	399 
    -- CP-element group 401:  members (9) 
      -- CP-element group 401: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Update/word_access_complete/word_0/ca
      -- CP-element group 401: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_update_completed_
      -- CP-element group 401: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Update/word_access_complete/word_0/$exit
      -- CP-element group 401: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Update/ptr_deref_798_Merge/merge_ack
      -- CP-element group 401: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Update/ptr_deref_798_Merge/$entry
      -- CP-element group 401: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Update/ptr_deref_798_Merge/$exit
      -- CP-element group 401: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Update/ptr_deref_798_Merge/merge_req
      -- CP-element group 401: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Update/$exit
      -- CP-element group 401: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_Update/word_access_complete/$exit
      -- 
    ca_1813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_798_load_0_ack_1, ack => zeropad_CP_182_elements(401)); -- 
    -- CP-element group 402:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	142 
    -- CP-element group 402: 	163 
    -- CP-element group 402: 	226 
    -- CP-element group 402: marked-predecessors 
    -- CP-element group 402: 	404 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	404 
    -- CP-element group 402:  members (3) 
      -- CP-element group 402: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_835_sample_start_
      -- CP-element group 402: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_835_Sample/req
      -- CP-element group 402: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_835_Sample/$entry
      -- 
    req_1826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(402), ack => W_ifx_xthen180_ifx_xthen191_taken_807_delayed_12_0_833_inst_req_0); -- 
    zeropad_cp_element_group_402: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_402"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(226) & zeropad_CP_182_elements(404);
      gj_zeropad_cp_element_group_402 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(402), clk => clk, reset => reset); --
    end block;
    -- CP-element group 403:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	115 
    -- CP-element group 403: marked-predecessors 
    -- CP-element group 403: 	405 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	405 
    -- CP-element group 403:  members (3) 
      -- CP-element group 403: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_835_update_start_
      -- CP-element group 403: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_835_Update/req
      -- CP-element group 403: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_835_Update/$entry
      -- 
    req_1831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(403), ack => W_ifx_xthen180_ifx_xthen191_taken_807_delayed_12_0_833_inst_req_1); -- 
    zeropad_cp_element_group_403: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_403"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(405);
      gj_zeropad_cp_element_group_403 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(403), clk => clk, reset => reset); --
    end block;
    -- CP-element group 404:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	402 
    -- CP-element group 404: successors 
    -- CP-element group 404: marked-successors 
    -- CP-element group 404: 	138 
    -- CP-element group 404: 	159 
    -- CP-element group 404: 	222 
    -- CP-element group 404: 	402 
    -- CP-element group 404:  members (3) 
      -- CP-element group 404: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_835_sample_completed_
      -- CP-element group 404: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_835_Sample/ack
      -- CP-element group 404: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_835_Sample/$exit
      -- 
    ack_1827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen180_ifx_xthen191_taken_807_delayed_12_0_833_inst_ack_0, ack => zeropad_CP_182_elements(404)); -- 
    -- CP-element group 405:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	403 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	611 
    -- CP-element group 405: marked-successors 
    -- CP-element group 405: 	326 
    -- CP-element group 405: 	403 
    -- CP-element group 405:  members (3) 
      -- CP-element group 405: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_835_Update/ack
      -- CP-element group 405: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_835_Update/$exit
      -- CP-element group 405: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_835_update_completed_
      -- 
    ack_1832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen180_ifx_xthen191_taken_807_delayed_12_0_833_inst_ack_1, ack => zeropad_CP_182_elements(405)); -- 
    -- CP-element group 406:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	142 
    -- CP-element group 406: 	163 
    -- CP-element group 406: 	226 
    -- CP-element group 406: 	331 
    -- CP-element group 406: marked-predecessors 
    -- CP-element group 406: 	408 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	408 
    -- CP-element group 406:  members (3) 
      -- CP-element group 406: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_842_start/req
      -- CP-element group 406: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_842_start/$entry
      -- CP-element group 406: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_842_sample_start_
      -- 
    req_1840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(406), ack => MUX_842_inst_req_0); -- 
    zeropad_cp_element_group_406: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_406"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(226) & zeropad_CP_182_elements(331) & zeropad_CP_182_elements(408);
      gj_zeropad_cp_element_group_406 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(406), clk => clk, reset => reset); --
    end block;
    -- CP-element group 407:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	115 
    -- CP-element group 407: marked-predecessors 
    -- CP-element group 407: 	409 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	409 
    -- CP-element group 407:  members (3) 
      -- CP-element group 407: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_842_complete/req
      -- CP-element group 407: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_842_complete/$entry
      -- CP-element group 407: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_842_update_start_
      -- 
    req_1845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(407), ack => MUX_842_inst_req_1); -- 
    zeropad_cp_element_group_407: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_407"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(409);
      gj_zeropad_cp_element_group_407 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(407), clk => clk, reset => reset); --
    end block;
    -- CP-element group 408:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	406 
    -- CP-element group 408: successors 
    -- CP-element group 408: marked-successors 
    -- CP-element group 408: 	138 
    -- CP-element group 408: 	159 
    -- CP-element group 408: 	222 
    -- CP-element group 408: 	327 
    -- CP-element group 408: 	406 
    -- CP-element group 408:  members (3) 
      -- CP-element group 408: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_842_start/ack
      -- CP-element group 408: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_842_start/$exit
      -- CP-element group 408: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_842_sample_completed_
      -- 
    ack_1841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_842_inst_ack_0, ack => zeropad_CP_182_elements(408)); -- 
    -- CP-element group 409:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	407 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	611 
    -- CP-element group 409: marked-successors 
    -- CP-element group 409: 	326 
    -- CP-element group 409: 	407 
    -- CP-element group 409:  members (3) 
      -- CP-element group 409: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_842_complete/ack
      -- CP-element group 409: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_842_complete/$exit
      -- CP-element group 409: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_842_update_completed_
      -- 
    ack_1846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_842_inst_ack_1, ack => zeropad_CP_182_elements(409)); -- 
    -- CP-element group 410:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	142 
    -- CP-element group 410: 	163 
    -- CP-element group 410: 	226 
    -- CP-element group 410: 	247 
    -- CP-element group 410: marked-predecessors 
    -- CP-element group 410: 	412 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	412 
    -- CP-element group 410:  members (3) 
      -- CP-element group 410: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_854_Sample/rr
      -- CP-element group 410: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_854_Sample/$entry
      -- CP-element group 410: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_854_sample_start_
      -- 
    rr_1854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(410), ack => type_cast_854_inst_req_0); -- 
    zeropad_cp_element_group_410: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_410"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(226) & zeropad_CP_182_elements(247) & zeropad_CP_182_elements(412);
      gj_zeropad_cp_element_group_410 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(410), clk => clk, reset => reset); --
    end block;
    -- CP-element group 411:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: marked-predecessors 
    -- CP-element group 411: 	413 
    -- CP-element group 411: 	444 
    -- CP-element group 411: 	448 
    -- CP-element group 411: 	452 
    -- CP-element group 411: 	456 
    -- CP-element group 411: 	488 
    -- CP-element group 411: 	492 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	413 
    -- CP-element group 411:  members (3) 
      -- CP-element group 411: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_854_Update/cr
      -- CP-element group 411: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_854_Update/$entry
      -- CP-element group 411: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_854_update_start_
      -- 
    cr_1859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(411), ack => type_cast_854_inst_req_1); -- 
    zeropad_cp_element_group_411: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_411"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(413) & zeropad_CP_182_elements(444) & zeropad_CP_182_elements(448) & zeropad_CP_182_elements(452) & zeropad_CP_182_elements(456) & zeropad_CP_182_elements(488) & zeropad_CP_182_elements(492);
      gj_zeropad_cp_element_group_411 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(411), clk => clk, reset => reset); --
    end block;
    -- CP-element group 412:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	410 
    -- CP-element group 412: successors 
    -- CP-element group 412: marked-successors 
    -- CP-element group 412: 	138 
    -- CP-element group 412: 	159 
    -- CP-element group 412: 	222 
    -- CP-element group 412: 	243 
    -- CP-element group 412: 	410 
    -- CP-element group 412:  members (3) 
      -- CP-element group 412: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_854_Sample/ra
      -- CP-element group 412: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_854_Sample/$exit
      -- CP-element group 412: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_854_sample_completed_
      -- 
    ra_1855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_854_inst_ack_0, ack => zeropad_CP_182_elements(412)); -- 
    -- CP-element group 413:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	411 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	442 
    -- CP-element group 413: 	446 
    -- CP-element group 413: 	450 
    -- CP-element group 413: 	454 
    -- CP-element group 413: 	486 
    -- CP-element group 413: 	490 
    -- CP-element group 413: marked-successors 
    -- CP-element group 413: 	411 
    -- CP-element group 413:  members (3) 
      -- CP-element group 413: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_854_Update/ca
      -- CP-element group 413: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_854_Update/$exit
      -- CP-element group 413: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_854_update_completed_
      -- 
    ca_1860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_854_inst_ack_1, ack => zeropad_CP_182_elements(413)); -- 
    -- CP-element group 414:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	142 
    -- CP-element group 414: 	163 
    -- CP-element group 414: 	226 
    -- CP-element group 414: marked-predecessors 
    -- CP-element group 414: 	416 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	416 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_858_Sample/req
      -- CP-element group 414: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_858_Sample/$entry
      -- CP-element group 414: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_858_sample_start_
      -- 
    req_1868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(414), ack => W_ifx_xthen191_exec_guard_823_delayed_1_0_856_inst_req_0); -- 
    zeropad_cp_element_group_414: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_414"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(226) & zeropad_CP_182_elements(416);
      gj_zeropad_cp_element_group_414 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(414), clk => clk, reset => reset); --
    end block;
    -- CP-element group 415:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: marked-predecessors 
    -- CP-element group 415: 	417 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	417 
    -- CP-element group 415:  members (3) 
      -- CP-element group 415: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_858_Update/req
      -- CP-element group 415: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_858_Update/$entry
      -- CP-element group 415: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_858_update_start_
      -- 
    req_1873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(415), ack => W_ifx_xthen191_exec_guard_823_delayed_1_0_856_inst_req_1); -- 
    zeropad_cp_element_group_415: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_415"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_CP_182_elements(417);
      gj_zeropad_cp_element_group_415 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(415), clk => clk, reset => reset); --
    end block;
    -- CP-element group 416:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	414 
    -- CP-element group 416: successors 
    -- CP-element group 416: marked-successors 
    -- CP-element group 416: 	138 
    -- CP-element group 416: 	159 
    -- CP-element group 416: 	222 
    -- CP-element group 416: 	414 
    -- CP-element group 416:  members (3) 
      -- CP-element group 416: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_858_Sample/ack
      -- CP-element group 416: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_858_Sample/$exit
      -- CP-element group 416: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_858_sample_completed_
      -- 
    ack_1869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen191_exec_guard_823_delayed_1_0_856_inst_ack_0, ack => zeropad_CP_182_elements(416)); -- 
    -- CP-element group 417:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	415 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	611 
    -- CP-element group 417: marked-successors 
    -- CP-element group 417: 	415 
    -- CP-element group 417:  members (3) 
      -- CP-element group 417: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_858_Update/$exit
      -- CP-element group 417: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_858_Update/ack
      -- CP-element group 417: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_858_update_completed_
      -- 
    ack_1874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen191_exec_guard_823_delayed_1_0_856_inst_ack_1, ack => zeropad_CP_182_elements(417)); -- 
    -- CP-element group 418:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	142 
    -- CP-element group 418: 	163 
    -- CP-element group 418: 	226 
    -- CP-element group 418: marked-predecessors 
    -- CP-element group 418: 	420 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	420 
    -- CP-element group 418:  members (3) 
      -- CP-element group 418: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_867_Sample/$entry
      -- CP-element group 418: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_867_sample_start_
      -- CP-element group 418: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_867_Sample/req
      -- 
    req_1882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(418), ack => W_ifx_xthen191_exec_guard_829_delayed_1_0_865_inst_req_0); -- 
    zeropad_cp_element_group_418: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_418"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(226) & zeropad_CP_182_elements(420);
      gj_zeropad_cp_element_group_418 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(418), clk => clk, reset => reset); --
    end block;
    -- CP-element group 419:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: marked-predecessors 
    -- CP-element group 419: 	421 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	421 
    -- CP-element group 419:  members (3) 
      -- CP-element group 419: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_867_Update/$entry
      -- CP-element group 419: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_867_update_start_
      -- CP-element group 419: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_867_Update/req
      -- 
    req_1887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(419), ack => W_ifx_xthen191_exec_guard_829_delayed_1_0_865_inst_req_1); -- 
    zeropad_cp_element_group_419: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_419"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_CP_182_elements(421);
      gj_zeropad_cp_element_group_419 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(419), clk => clk, reset => reset); --
    end block;
    -- CP-element group 420:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	418 
    -- CP-element group 420: successors 
    -- CP-element group 420: marked-successors 
    -- CP-element group 420: 	138 
    -- CP-element group 420: 	159 
    -- CP-element group 420: 	222 
    -- CP-element group 420: 	418 
    -- CP-element group 420:  members (3) 
      -- CP-element group 420: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_867_Sample/ack
      -- CP-element group 420: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_867_sample_completed_
      -- CP-element group 420: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_867_Sample/$exit
      -- 
    ack_1883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen191_exec_guard_829_delayed_1_0_865_inst_ack_0, ack => zeropad_CP_182_elements(420)); -- 
    -- CP-element group 421:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	419 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	611 
    -- CP-element group 421: marked-successors 
    -- CP-element group 421: 	419 
    -- CP-element group 421:  members (3) 
      -- CP-element group 421: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_867_update_completed_
      -- CP-element group 421: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_867_Update/$exit
      -- CP-element group 421: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_867_Update/ack
      -- 
    ack_1888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen191_exec_guard_829_delayed_1_0_865_inst_ack_1, ack => zeropad_CP_182_elements(421)); -- 
    -- CP-element group 422:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	112 
    -- CP-element group 422: marked-predecessors 
    -- CP-element group 422: 	424 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	424 
    -- CP-element group 422:  members (3) 
      -- CP-element group 422: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_871_Sample/$entry
      -- CP-element group 422: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_871_sample_start_
      -- CP-element group 422: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_871_Sample/rr
      -- 
    rr_1896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(422), ack => type_cast_871_inst_req_0); -- 
    zeropad_cp_element_group_422: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_422"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(424);
      gj_zeropad_cp_element_group_422 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(422), clk => clk, reset => reset); --
    end block;
    -- CP-element group 423:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: marked-predecessors 
    -- CP-element group 423: 	425 
    -- CP-element group 423: 	444 
    -- CP-element group 423: 	448 
    -- CP-element group 423: 	452 
    -- CP-element group 423: 	456 
    -- CP-element group 423: 	488 
    -- CP-element group 423: 	492 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	425 
    -- CP-element group 423:  members (3) 
      -- CP-element group 423: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_871_update_start_
      -- CP-element group 423: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_871_Update/$entry
      -- CP-element group 423: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_871_Update/cr
      -- 
    cr_1901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(423), ack => type_cast_871_inst_req_1); -- 
    zeropad_cp_element_group_423: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_423"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(425) & zeropad_CP_182_elements(444) & zeropad_CP_182_elements(448) & zeropad_CP_182_elements(452) & zeropad_CP_182_elements(456) & zeropad_CP_182_elements(488) & zeropad_CP_182_elements(492);
      gj_zeropad_cp_element_group_423 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(423), clk => clk, reset => reset); --
    end block;
    -- CP-element group 424:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	422 
    -- CP-element group 424: successors 
    -- CP-element group 424: marked-successors 
    -- CP-element group 424: 	422 
    -- CP-element group 424:  members (3) 
      -- CP-element group 424: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_871_Sample/ra
      -- CP-element group 424: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_871_Sample/$exit
      -- CP-element group 424: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_871_sample_completed_
      -- 
    ra_1897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_871_inst_ack_0, ack => zeropad_CP_182_elements(424)); -- 
    -- CP-element group 425:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	423 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	442 
    -- CP-element group 425: 	446 
    -- CP-element group 425: 	450 
    -- CP-element group 425: 	454 
    -- CP-element group 425: 	486 
    -- CP-element group 425: 	490 
    -- CP-element group 425: marked-successors 
    -- CP-element group 425: 	423 
    -- CP-element group 425:  members (3) 
      -- CP-element group 425: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_871_Update/ca
      -- CP-element group 425: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_871_update_completed_
      -- CP-element group 425: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_871_Update/$exit
      -- 
    ca_1902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 425_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_871_inst_ack_1, ack => zeropad_CP_182_elements(425)); -- 
    -- CP-element group 426:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	142 
    -- CP-element group 426: 	163 
    -- CP-element group 426: 	226 
    -- CP-element group 426: marked-predecessors 
    -- CP-element group 426: 	428 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	428 
    -- CP-element group 426:  members (3) 
      -- CP-element group 426: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_882_sample_start_
      -- CP-element group 426: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_882_Sample/$entry
      -- CP-element group 426: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_882_Sample/req
      -- 
    req_1910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(426), ack => W_ifx_xthen191_exec_guard_838_delayed_1_0_880_inst_req_0); -- 
    zeropad_cp_element_group_426: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_426"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(226) & zeropad_CP_182_elements(428);
      gj_zeropad_cp_element_group_426 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(426), clk => clk, reset => reset); --
    end block;
    -- CP-element group 427:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: marked-predecessors 
    -- CP-element group 427: 	429 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	429 
    -- CP-element group 427:  members (3) 
      -- CP-element group 427: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_882_update_start_
      -- CP-element group 427: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_882_Update/$entry
      -- CP-element group 427: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_882_Update/req
      -- 
    req_1915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(427), ack => W_ifx_xthen191_exec_guard_838_delayed_1_0_880_inst_req_1); -- 
    zeropad_cp_element_group_427: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_427"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_CP_182_elements(429);
      gj_zeropad_cp_element_group_427 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(427), clk => clk, reset => reset); --
    end block;
    -- CP-element group 428:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	426 
    -- CP-element group 428: successors 
    -- CP-element group 428: marked-successors 
    -- CP-element group 428: 	138 
    -- CP-element group 428: 	159 
    -- CP-element group 428: 	222 
    -- CP-element group 428: 	426 
    -- CP-element group 428:  members (3) 
      -- CP-element group 428: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_882_sample_completed_
      -- CP-element group 428: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_882_Sample/$exit
      -- CP-element group 428: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_882_Sample/ack
      -- 
    ack_1911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen191_exec_guard_838_delayed_1_0_880_inst_ack_0, ack => zeropad_CP_182_elements(428)); -- 
    -- CP-element group 429:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	427 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	611 
    -- CP-element group 429: marked-successors 
    -- CP-element group 429: 	427 
    -- CP-element group 429:  members (3) 
      -- CP-element group 429: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_882_update_completed_
      -- CP-element group 429: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_882_Update/$exit
      -- CP-element group 429: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_882_Update/ack
      -- 
    ack_1916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 429_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen191_exec_guard_838_delayed_1_0_880_inst_ack_1, ack => zeropad_CP_182_elements(429)); -- 
    -- CP-element group 430:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	142 
    -- CP-element group 430: 	163 
    -- CP-element group 430: 	226 
    -- CP-element group 430: marked-predecessors 
    -- CP-element group 430: 	432 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	432 
    -- CP-element group 430:  members (3) 
      -- CP-element group 430: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_891_sample_start_
      -- CP-element group 430: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_891_Sample/$entry
      -- CP-element group 430: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_891_Sample/req
      -- 
    req_1924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(430), ack => W_ifx_xthen191_exec_guard_845_delayed_1_0_889_inst_req_0); -- 
    zeropad_cp_element_group_430: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_430"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(226) & zeropad_CP_182_elements(432);
      gj_zeropad_cp_element_group_430 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(430), clk => clk, reset => reset); --
    end block;
    -- CP-element group 431:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: marked-predecessors 
    -- CP-element group 431: 	433 
    -- CP-element group 431: 	488 
    -- CP-element group 431: 	492 
    -- CP-element group 431: successors 
    -- CP-element group 431: 	433 
    -- CP-element group 431:  members (3) 
      -- CP-element group 431: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_891_update_start_
      -- CP-element group 431: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_891_Update/$entry
      -- CP-element group 431: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_891_Update/req
      -- 
    req_1929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(431), ack => W_ifx_xthen191_exec_guard_845_delayed_1_0_889_inst_req_1); -- 
    zeropad_cp_element_group_431: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_431"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(433) & zeropad_CP_182_elements(488) & zeropad_CP_182_elements(492);
      gj_zeropad_cp_element_group_431 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(431), clk => clk, reset => reset); --
    end block;
    -- CP-element group 432:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	430 
    -- CP-element group 432: successors 
    -- CP-element group 432: marked-successors 
    -- CP-element group 432: 	138 
    -- CP-element group 432: 	159 
    -- CP-element group 432: 	222 
    -- CP-element group 432: 	430 
    -- CP-element group 432:  members (3) 
      -- CP-element group 432: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_891_Sample/$exit
      -- CP-element group 432: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_891_sample_completed_
      -- CP-element group 432: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_891_Sample/ack
      -- 
    ack_1925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen191_exec_guard_845_delayed_1_0_889_inst_ack_0, ack => zeropad_CP_182_elements(432)); -- 
    -- CP-element group 433:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	431 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	486 
    -- CP-element group 433: 	490 
    -- CP-element group 433: marked-successors 
    -- CP-element group 433: 	431 
    -- CP-element group 433:  members (3) 
      -- CP-element group 433: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_891_update_completed_
      -- CP-element group 433: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_891_Update/$exit
      -- CP-element group 433: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_891_Update/ack
      -- 
    ack_1930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 433_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen191_exec_guard_845_delayed_1_0_889_inst_ack_1, ack => zeropad_CP_182_elements(433)); -- 
    -- CP-element group 434:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	142 
    -- CP-element group 434: 	163 
    -- CP-element group 434: 	226 
    -- CP-element group 434: marked-predecessors 
    -- CP-element group 434: 	436 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	436 
    -- CP-element group 434:  members (3) 
      -- CP-element group 434: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_899_Sample/req
      -- CP-element group 434: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_899_sample_start_
      -- CP-element group 434: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_899_Sample/$entry
      -- 
    req_1938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(434), ack => W_ifx_xthen191_exec_guard_850_delayed_1_0_897_inst_req_0); -- 
    zeropad_cp_element_group_434: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_434"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(226) & zeropad_CP_182_elements(436);
      gj_zeropad_cp_element_group_434 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(434), clk => clk, reset => reset); --
    end block;
    -- CP-element group 435:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: marked-predecessors 
    -- CP-element group 435: 	437 
    -- CP-element group 435: 	444 
    -- CP-element group 435: 	448 
    -- CP-element group 435: 	452 
    -- CP-element group 435: 	456 
    -- CP-element group 435: successors 
    -- CP-element group 435: 	437 
    -- CP-element group 435:  members (3) 
      -- CP-element group 435: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_899_Update/req
      -- CP-element group 435: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_899_Update/$entry
      -- CP-element group 435: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_899_update_start_
      -- 
    req_1943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(435), ack => W_ifx_xthen191_exec_guard_850_delayed_1_0_897_inst_req_1); -- 
    zeropad_cp_element_group_435: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_435"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(437) & zeropad_CP_182_elements(444) & zeropad_CP_182_elements(448) & zeropad_CP_182_elements(452) & zeropad_CP_182_elements(456);
      gj_zeropad_cp_element_group_435 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(435), clk => clk, reset => reset); --
    end block;
    -- CP-element group 436:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	434 
    -- CP-element group 436: successors 
    -- CP-element group 436: marked-successors 
    -- CP-element group 436: 	138 
    -- CP-element group 436: 	159 
    -- CP-element group 436: 	222 
    -- CP-element group 436: 	434 
    -- CP-element group 436:  members (3) 
      -- CP-element group 436: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_899_Sample/ack
      -- CP-element group 436: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_899_sample_completed_
      -- CP-element group 436: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_899_Sample/$exit
      -- 
    ack_1939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen191_exec_guard_850_delayed_1_0_897_inst_ack_0, ack => zeropad_CP_182_elements(436)); -- 
    -- CP-element group 437:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	435 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	442 
    -- CP-element group 437: 	446 
    -- CP-element group 437: 	450 
    -- CP-element group 437: 	454 
    -- CP-element group 437: marked-successors 
    -- CP-element group 437: 	435 
    -- CP-element group 437:  members (3) 
      -- CP-element group 437: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_899_Update/$exit
      -- CP-element group 437: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_899_Update/ack
      -- CP-element group 437: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_899_update_completed_
      -- 
    ack_1944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 437_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen191_exec_guard_850_delayed_1_0_897_inst_ack_1, ack => zeropad_CP_182_elements(437)); -- 
    -- CP-element group 438:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	268 
    -- CP-element group 438: marked-predecessors 
    -- CP-element group 438: 	440 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	440 
    -- CP-element group 438:  members (3) 
      -- CP-element group 438: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_911_Sample/req
      -- CP-element group 438: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_911_sample_start_
      -- CP-element group 438: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_911_Sample/$entry
      -- 
    req_1952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(438), ack => W_o1x_x1_860_delayed_1_0_909_inst_req_0); -- 
    zeropad_cp_element_group_438: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_438"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(268) & zeropad_CP_182_elements(440);
      gj_zeropad_cp_element_group_438 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(438), clk => clk, reset => reset); --
    end block;
    -- CP-element group 439:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: marked-predecessors 
    -- CP-element group 439: 	441 
    -- CP-element group 439: 	444 
    -- CP-element group 439: successors 
    -- CP-element group 439: 	441 
    -- CP-element group 439:  members (3) 
      -- CP-element group 439: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_911_update_start_
      -- CP-element group 439: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_911_Update/$entry
      -- CP-element group 439: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_911_Update/req
      -- 
    req_1957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(439), ack => W_o1x_x1_860_delayed_1_0_909_inst_req_1); -- 
    zeropad_cp_element_group_439: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_439"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(441) & zeropad_CP_182_elements(444);
      gj_zeropad_cp_element_group_439 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(439), clk => clk, reset => reset); --
    end block;
    -- CP-element group 440:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	438 
    -- CP-element group 440: successors 
    -- CP-element group 440: marked-successors 
    -- CP-element group 440: 	264 
    -- CP-element group 440: 	438 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_911_Sample/ack
      -- CP-element group 440: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_911_sample_completed_
      -- CP-element group 440: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_911_Sample/$exit
      -- 
    ack_1953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_o1x_x1_860_delayed_1_0_909_inst_ack_0, ack => zeropad_CP_182_elements(440)); -- 
    -- CP-element group 441:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	439 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	442 
    -- CP-element group 441: marked-successors 
    -- CP-element group 441: 	439 
    -- CP-element group 441:  members (3) 
      -- CP-element group 441: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_911_update_completed_
      -- CP-element group 441: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_911_Update/$exit
      -- CP-element group 441: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_911_Update/ack
      -- 
    ack_1958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 441_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_o1x_x1_860_delayed_1_0_909_inst_ack_1, ack => zeropad_CP_182_elements(441)); -- 
    -- CP-element group 442:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	413 
    -- CP-element group 442: 	425 
    -- CP-element group 442: 	437 
    -- CP-element group 442: 	441 
    -- CP-element group 442: marked-predecessors 
    -- CP-element group 442: 	444 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	444 
    -- CP-element group 442:  members (3) 
      -- CP-element group 442: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_915_Sample/$entry
      -- CP-element group 442: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_915_Sample/rr
      -- CP-element group 442: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_915_sample_start_
      -- 
    rr_1966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(442), ack => type_cast_915_inst_req_0); -- 
    zeropad_cp_element_group_442: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_442"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(413) & zeropad_CP_182_elements(425) & zeropad_CP_182_elements(437) & zeropad_CP_182_elements(441) & zeropad_CP_182_elements(444);
      gj_zeropad_cp_element_group_442 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(442), clk => clk, reset => reset); --
    end block;
    -- CP-element group 443:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	115 
    -- CP-element group 443: marked-predecessors 
    -- CP-element group 443: 	445 
    -- CP-element group 443: 	464 
    -- CP-element group 443: 	472 
    -- CP-element group 443: 	476 
    -- CP-element group 443: 	500 
    -- CP-element group 443: 	508 
    -- CP-element group 443: 	512 
    -- CP-element group 443: 	520 
    -- CP-element group 443: 	548 
    -- CP-element group 443: 	571 
    -- CP-element group 443: successors 
    -- CP-element group 443: 	445 
    -- CP-element group 443:  members (3) 
      -- CP-element group 443: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_915_Update/cr
      -- CP-element group 443: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_915_update_start_
      -- CP-element group 443: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_915_Update/$entry
      -- 
    cr_1971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(443), ack => type_cast_915_inst_req_1); -- 
    zeropad_cp_element_group_443: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_443"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(445) & zeropad_CP_182_elements(464) & zeropad_CP_182_elements(472) & zeropad_CP_182_elements(476) & zeropad_CP_182_elements(500) & zeropad_CP_182_elements(508) & zeropad_CP_182_elements(512) & zeropad_CP_182_elements(520) & zeropad_CP_182_elements(548) & zeropad_CP_182_elements(571);
      gj_zeropad_cp_element_group_443 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(443), clk => clk, reset => reset); --
    end block;
    -- CP-element group 444:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	442 
    -- CP-element group 444: successors 
    -- CP-element group 444: marked-successors 
    -- CP-element group 444: 	411 
    -- CP-element group 444: 	423 
    -- CP-element group 444: 	435 
    -- CP-element group 444: 	439 
    -- CP-element group 444: 	442 
    -- CP-element group 444:  members (3) 
      -- CP-element group 444: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_915_sample_completed_
      -- CP-element group 444: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_915_Sample/$exit
      -- CP-element group 444: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_915_Sample/ra
      -- 
    ra_1967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_915_inst_ack_0, ack => zeropad_CP_182_elements(444)); -- 
    -- CP-element group 445:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	443 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	462 
    -- CP-element group 445: 	470 
    -- CP-element group 445: 	474 
    -- CP-element group 445: 	498 
    -- CP-element group 445: 	506 
    -- CP-element group 445: 	510 
    -- CP-element group 445: 	518 
    -- CP-element group 445: 	546 
    -- CP-element group 445: 	569 
    -- CP-element group 445: marked-successors 
    -- CP-element group 445: 	118 
    -- CP-element group 445: 	179 
    -- CP-element group 445: 	200 
    -- CP-element group 445: 	221 
    -- CP-element group 445: 	305 
    -- CP-element group 445: 	443 
    -- CP-element group 445:  members (3) 
      -- CP-element group 445: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_915_Update/$exit
      -- CP-element group 445: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_915_Update/ca
      -- CP-element group 445: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_915_update_completed_
      -- 
    ca_1972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 445_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_915_inst_ack_1, ack => zeropad_CP_182_elements(445)); -- 
    -- CP-element group 446:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	413 
    -- CP-element group 446: 	425 
    -- CP-element group 446: 	437 
    -- CP-element group 446: marked-predecessors 
    -- CP-element group 446: 	448 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	448 
    -- CP-element group 446:  members (3) 
      -- CP-element group 446: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_919_Sample/req
      -- CP-element group 446: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_919_Sample/$entry
      -- CP-element group 446: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_919_sample_start_
      -- 
    req_1980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(446), ack => W_landx_xlhsx_xtrue208_exec_guard_863_delayed_1_0_917_inst_req_0); -- 
    zeropad_cp_element_group_446: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_446"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(413) & zeropad_CP_182_elements(425) & zeropad_CP_182_elements(437) & zeropad_CP_182_elements(448);
      gj_zeropad_cp_element_group_446 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(446), clk => clk, reset => reset); --
    end block;
    -- CP-element group 447:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: marked-predecessors 
    -- CP-element group 447: 	449 
    -- CP-element group 447: successors 
    -- CP-element group 447: 	449 
    -- CP-element group 447:  members (3) 
      -- CP-element group 447: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_919_Update/req
      -- CP-element group 447: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_919_Update/$entry
      -- CP-element group 447: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_919_update_start_
      -- 
    req_1985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(447), ack => W_landx_xlhsx_xtrue208_exec_guard_863_delayed_1_0_917_inst_req_1); -- 
    zeropad_cp_element_group_447: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_447"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_CP_182_elements(449);
      gj_zeropad_cp_element_group_447 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(447), clk => clk, reset => reset); --
    end block;
    -- CP-element group 448:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	446 
    -- CP-element group 448: successors 
    -- CP-element group 448: marked-successors 
    -- CP-element group 448: 	411 
    -- CP-element group 448: 	423 
    -- CP-element group 448: 	435 
    -- CP-element group 448: 	446 
    -- CP-element group 448:  members (3) 
      -- CP-element group 448: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_919_Sample/ack
      -- CP-element group 448: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_919_Sample/$exit
      -- CP-element group 448: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_919_sample_completed_
      -- 
    ack_1981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 448_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue208_exec_guard_863_delayed_1_0_917_inst_ack_0, ack => zeropad_CP_182_elements(448)); -- 
    -- CP-element group 449:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	447 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	611 
    -- CP-element group 449: marked-successors 
    -- CP-element group 449: 	447 
    -- CP-element group 449:  members (3) 
      -- CP-element group 449: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_919_Update/ack
      -- CP-element group 449: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_919_Update/$exit
      -- CP-element group 449: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_919_update_completed_
      -- 
    ack_1986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 449_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue208_exec_guard_863_delayed_1_0_917_inst_ack_1, ack => zeropad_CP_182_elements(449)); -- 
    -- CP-element group 450:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	413 
    -- CP-element group 450: 	425 
    -- CP-element group 450: 	437 
    -- CP-element group 450: marked-predecessors 
    -- CP-element group 450: 	452 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	452 
    -- CP-element group 450:  members (3) 
      -- CP-element group 450: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_928_sample_start_
      -- CP-element group 450: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_928_Sample/$entry
      -- CP-element group 450: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_928_Sample/req
      -- 
    req_1994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(450), ack => W_landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_926_inst_req_0); -- 
    zeropad_cp_element_group_450: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_450"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(413) & zeropad_CP_182_elements(425) & zeropad_CP_182_elements(437) & zeropad_CP_182_elements(452);
      gj_zeropad_cp_element_group_450 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(450), clk => clk, reset => reset); --
    end block;
    -- CP-element group 451:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	115 
    -- CP-element group 451: marked-predecessors 
    -- CP-element group 451: 	453 
    -- CP-element group 451: 	464 
    -- CP-element group 451: 	472 
    -- CP-element group 451: 	476 
    -- CP-element group 451: 	508 
    -- CP-element group 451: 	512 
    -- CP-element group 451: 	520 
    -- CP-element group 451: 	548 
    -- CP-element group 451: 	571 
    -- CP-element group 451: successors 
    -- CP-element group 451: 	453 
    -- CP-element group 451:  members (3) 
      -- CP-element group 451: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_928_update_start_
      -- CP-element group 451: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_928_Update/$entry
      -- CP-element group 451: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_928_Update/req
      -- 
    req_1999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(451), ack => W_landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_926_inst_req_1); -- 
    zeropad_cp_element_group_451: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_451"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(453) & zeropad_CP_182_elements(464) & zeropad_CP_182_elements(472) & zeropad_CP_182_elements(476) & zeropad_CP_182_elements(508) & zeropad_CP_182_elements(512) & zeropad_CP_182_elements(520) & zeropad_CP_182_elements(548) & zeropad_CP_182_elements(571);
      gj_zeropad_cp_element_group_451 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(451), clk => clk, reset => reset); --
    end block;
    -- CP-element group 452:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	450 
    -- CP-element group 452: successors 
    -- CP-element group 452: marked-successors 
    -- CP-element group 452: 	411 
    -- CP-element group 452: 	423 
    -- CP-element group 452: 	435 
    -- CP-element group 452: 	450 
    -- CP-element group 452:  members (3) 
      -- CP-element group 452: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_928_sample_completed_
      -- CP-element group 452: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_928_Sample/$exit
      -- CP-element group 452: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_928_Sample/ack
      -- 
    ack_1995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 452_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_926_inst_ack_0, ack => zeropad_CP_182_elements(452)); -- 
    -- CP-element group 453:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	451 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	462 
    -- CP-element group 453: 	470 
    -- CP-element group 453: 	474 
    -- CP-element group 453: 	506 
    -- CP-element group 453: 	510 
    -- CP-element group 453: 	518 
    -- CP-element group 453: 	546 
    -- CP-element group 453: 	569 
    -- CP-element group 453: marked-successors 
    -- CP-element group 453: 	118 
    -- CP-element group 453: 	179 
    -- CP-element group 453: 	200 
    -- CP-element group 453: 	221 
    -- CP-element group 453: 	305 
    -- CP-element group 453: 	451 
    -- CP-element group 453:  members (3) 
      -- CP-element group 453: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_928_update_completed_
      -- CP-element group 453: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_928_Update/$exit
      -- CP-element group 453: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_928_Update/ack
      -- 
    ack_2000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 453_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_926_inst_ack_1, ack => zeropad_CP_182_elements(453)); -- 
    -- CP-element group 454:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	413 
    -- CP-element group 454: 	425 
    -- CP-element group 454: 	437 
    -- CP-element group 454: marked-predecessors 
    -- CP-element group 454: 	456 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	456 
    -- CP-element group 454:  members (3) 
      -- CP-element group 454: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_936_sample_start_
      -- CP-element group 454: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_936_Sample/$entry
      -- CP-element group 454: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_936_Sample/req
      -- 
    req_2008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(454), ack => W_landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_934_inst_req_0); -- 
    zeropad_cp_element_group_454: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_454"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(413) & zeropad_CP_182_elements(425) & zeropad_CP_182_elements(437) & zeropad_CP_182_elements(456);
      gj_zeropad_cp_element_group_454 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(454), clk => clk, reset => reset); --
    end block;
    -- CP-element group 455:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	115 
    -- CP-element group 455: marked-predecessors 
    -- CP-element group 455: 	457 
    -- CP-element group 455: 	500 
    -- CP-element group 455: 	512 
    -- CP-element group 455: 	520 
    -- CP-element group 455: 	548 
    -- CP-element group 455: 	571 
    -- CP-element group 455: successors 
    -- CP-element group 455: 	457 
    -- CP-element group 455:  members (3) 
      -- CP-element group 455: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_936_update_start_
      -- CP-element group 455: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_936_Update/$entry
      -- CP-element group 455: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_936_Update/req
      -- 
    req_2013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(455), ack => W_landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_934_inst_req_1); -- 
    zeropad_cp_element_group_455: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_455"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(457) & zeropad_CP_182_elements(500) & zeropad_CP_182_elements(512) & zeropad_CP_182_elements(520) & zeropad_CP_182_elements(548) & zeropad_CP_182_elements(571);
      gj_zeropad_cp_element_group_455 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(455), clk => clk, reset => reset); --
    end block;
    -- CP-element group 456:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	454 
    -- CP-element group 456: successors 
    -- CP-element group 456: marked-successors 
    -- CP-element group 456: 	411 
    -- CP-element group 456: 	423 
    -- CP-element group 456: 	435 
    -- CP-element group 456: 	454 
    -- CP-element group 456:  members (3) 
      -- CP-element group 456: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_936_sample_completed_
      -- CP-element group 456: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_936_Sample/$exit
      -- CP-element group 456: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_936_Sample/ack
      -- 
    ack_2009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 456_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_934_inst_ack_0, ack => zeropad_CP_182_elements(456)); -- 
    -- CP-element group 457:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	455 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	498 
    -- CP-element group 457: 	510 
    -- CP-element group 457: 	518 
    -- CP-element group 457: 	546 
    -- CP-element group 457: 	569 
    -- CP-element group 457: marked-successors 
    -- CP-element group 457: 	118 
    -- CP-element group 457: 	179 
    -- CP-element group 457: 	200 
    -- CP-element group 457: 	221 
    -- CP-element group 457: 	305 
    -- CP-element group 457: 	455 
    -- CP-element group 457:  members (3) 
      -- CP-element group 457: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_936_update_completed_
      -- CP-element group 457: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_936_Update/$exit
      -- CP-element group 457: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_936_Update/ack
      -- 
    ack_2014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 457_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_934_inst_ack_1, ack => zeropad_CP_182_elements(457)); -- 
    -- CP-element group 458:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	289 
    -- CP-element group 458: marked-predecessors 
    -- CP-element group 458: 	460 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	460 
    -- CP-element group 458:  members (3) 
      -- CP-element group 458: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_948_sample_start_
      -- CP-element group 458: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_948_Sample/$entry
      -- CP-element group 458: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_948_Sample/req
      -- 
    req_2022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(458), ack => W_o2x_x1_885_delayed_2_0_946_inst_req_0); -- 
    zeropad_cp_element_group_458: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_458"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(289) & zeropad_CP_182_elements(460);
      gj_zeropad_cp_element_group_458 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(458), clk => clk, reset => reset); --
    end block;
    -- CP-element group 459:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: marked-predecessors 
    -- CP-element group 459: 	461 
    -- CP-element group 459: 	464 
    -- CP-element group 459: successors 
    -- CP-element group 459: 	461 
    -- CP-element group 459:  members (3) 
      -- CP-element group 459: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_948_update_start_
      -- CP-element group 459: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_948_Update/$entry
      -- CP-element group 459: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_948_Update/req
      -- 
    req_2027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(459), ack => W_o2x_x1_885_delayed_2_0_946_inst_req_1); -- 
    zeropad_cp_element_group_459: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_459"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(461) & zeropad_CP_182_elements(464);
      gj_zeropad_cp_element_group_459 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(459), clk => clk, reset => reset); --
    end block;
    -- CP-element group 460:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	458 
    -- CP-element group 460: successors 
    -- CP-element group 460: marked-successors 
    -- CP-element group 460: 	285 
    -- CP-element group 460: 	458 
    -- CP-element group 460:  members (3) 
      -- CP-element group 460: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_948_sample_completed_
      -- CP-element group 460: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_948_Sample/$exit
      -- CP-element group 460: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_948_Sample/ack
      -- 
    ack_2023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 460_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_o2x_x1_885_delayed_2_0_946_inst_ack_0, ack => zeropad_CP_182_elements(460)); -- 
    -- CP-element group 461:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	459 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	462 
    -- CP-element group 461: marked-successors 
    -- CP-element group 461: 	459 
    -- CP-element group 461:  members (3) 
      -- CP-element group 461: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_948_update_completed_
      -- CP-element group 461: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_948_Update/$exit
      -- CP-element group 461: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_948_Update/ack
      -- 
    ack_2028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 461_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_o2x_x1_885_delayed_2_0_946_inst_ack_1, ack => zeropad_CP_182_elements(461)); -- 
    -- CP-element group 462:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	445 
    -- CP-element group 462: 	453 
    -- CP-element group 462: 	461 
    -- CP-element group 462: marked-predecessors 
    -- CP-element group 462: 	464 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	464 
    -- CP-element group 462:  members (3) 
      -- CP-element group 462: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_952_sample_start_
      -- CP-element group 462: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_952_Sample/$entry
      -- CP-element group 462: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_952_Sample/rr
      -- 
    rr_2036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(462), ack => type_cast_952_inst_req_0); -- 
    zeropad_cp_element_group_462: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_462"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(445) & zeropad_CP_182_elements(453) & zeropad_CP_182_elements(461) & zeropad_CP_182_elements(464);
      gj_zeropad_cp_element_group_462 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(462), clk => clk, reset => reset); --
    end block;
    -- CP-element group 463:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	115 
    -- CP-element group 463: marked-predecessors 
    -- CP-element group 463: 	465 
    -- CP-element group 463: successors 
    -- CP-element group 463: 	465 
    -- CP-element group 463:  members (3) 
      -- CP-element group 463: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_952_update_start_
      -- CP-element group 463: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_952_Update/$entry
      -- CP-element group 463: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_952_Update/cr
      -- 
    cr_2041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(463), ack => type_cast_952_inst_req_1); -- 
    zeropad_cp_element_group_463: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_463"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(465);
      gj_zeropad_cp_element_group_463 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(463), clk => clk, reset => reset); --
    end block;
    -- CP-element group 464:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	462 
    -- CP-element group 464: successors 
    -- CP-element group 464: marked-successors 
    -- CP-element group 464: 	443 
    -- CP-element group 464: 	451 
    -- CP-element group 464: 	459 
    -- CP-element group 464: 	462 
    -- CP-element group 464:  members (3) 
      -- CP-element group 464: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_952_sample_completed_
      -- CP-element group 464: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_952_Sample/$exit
      -- CP-element group 464: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_952_Sample/ra
      -- 
    ra_2037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 464_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_952_inst_ack_0, ack => zeropad_CP_182_elements(464)); -- 
    -- CP-element group 465:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	463 
    -- CP-element group 465: successors 
    -- CP-element group 465: 	611 
    -- CP-element group 465: marked-successors 
    -- CP-element group 465: 	137 
    -- CP-element group 465: 	463 
    -- CP-element group 465:  members (3) 
      -- CP-element group 465: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_952_update_completed_
      -- CP-element group 465: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_952_Update/$exit
      -- CP-element group 465: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_952_Update/ca
      -- 
    ca_2042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 465_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_952_inst_ack_1, ack => zeropad_CP_182_elements(465)); -- 
    -- CP-element group 466:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	142 
    -- CP-element group 466: marked-predecessors 
    -- CP-element group 466: 	468 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	468 
    -- CP-element group 466:  members (3) 
      -- CP-element group 466: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_956_sample_start_
      -- CP-element group 466: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_956_Sample/$entry
      -- CP-element group 466: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_956_Sample/req
      -- 
    req_2050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(466), ack => W_target_out_offsetx_x1_890_delayed_2_0_954_inst_req_0); -- 
    zeropad_cp_element_group_466: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_466"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(468);
      gj_zeropad_cp_element_group_466 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(466), clk => clk, reset => reset); --
    end block;
    -- CP-element group 467:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: marked-predecessors 
    -- CP-element group 467: 	469 
    -- CP-element group 467: 	480 
    -- CP-element group 467: successors 
    -- CP-element group 467: 	469 
    -- CP-element group 467:  members (3) 
      -- CP-element group 467: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_956_update_start_
      -- CP-element group 467: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_956_Update/$entry
      -- CP-element group 467: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_956_Update/req
      -- 
    req_2055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(467), ack => W_target_out_offsetx_x1_890_delayed_2_0_954_inst_req_1); -- 
    zeropad_cp_element_group_467: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_467"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(469) & zeropad_CP_182_elements(480);
      gj_zeropad_cp_element_group_467 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(467), clk => clk, reset => reset); --
    end block;
    -- CP-element group 468:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	466 
    -- CP-element group 468: successors 
    -- CP-element group 468: marked-successors 
    -- CP-element group 468: 	138 
    -- CP-element group 468: 	466 
    -- CP-element group 468:  members (3) 
      -- CP-element group 468: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_956_sample_completed_
      -- CP-element group 468: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_956_Sample/$exit
      -- CP-element group 468: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_956_Sample/ack
      -- 
    ack_2051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_target_out_offsetx_x1_890_delayed_2_0_954_inst_ack_0, ack => zeropad_CP_182_elements(468)); -- 
    -- CP-element group 469:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	467 
    -- CP-element group 469: successors 
    -- CP-element group 469: 	478 
    -- CP-element group 469: marked-successors 
    -- CP-element group 469: 	467 
    -- CP-element group 469:  members (3) 
      -- CP-element group 469: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_956_update_completed_
      -- CP-element group 469: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_956_Update/$exit
      -- CP-element group 469: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_956_Update/ack
      -- 
    ack_2056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 469_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_target_out_offsetx_x1_890_delayed_2_0_954_inst_ack_1, ack => zeropad_CP_182_elements(469)); -- 
    -- CP-element group 470:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	445 
    -- CP-element group 470: 	453 
    -- CP-element group 470: marked-predecessors 
    -- CP-element group 470: 	472 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	472 
    -- CP-element group 470:  members (3) 
      -- CP-element group 470: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_965_sample_start_
      -- CP-element group 470: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_965_Sample/$entry
      -- CP-element group 470: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_965_Sample/req
      -- 
    req_2064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(470), ack => W_landx_xlhsx_xtrue219_exec_guard_894_delayed_1_0_963_inst_req_0); -- 
    zeropad_cp_element_group_470: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_470"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(445) & zeropad_CP_182_elements(453) & zeropad_CP_182_elements(472);
      gj_zeropad_cp_element_group_470 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(470), clk => clk, reset => reset); --
    end block;
    -- CP-element group 471:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: marked-predecessors 
    -- CP-element group 471: 	473 
    -- CP-element group 471: successors 
    -- CP-element group 471: 	473 
    -- CP-element group 471:  members (3) 
      -- CP-element group 471: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_965_update_start_
      -- CP-element group 471: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_965_Update/$entry
      -- CP-element group 471: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_965_Update/req
      -- 
    req_2069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(471), ack => W_landx_xlhsx_xtrue219_exec_guard_894_delayed_1_0_963_inst_req_1); -- 
    zeropad_cp_element_group_471: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_471"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_CP_182_elements(473);
      gj_zeropad_cp_element_group_471 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(471), clk => clk, reset => reset); --
    end block;
    -- CP-element group 472:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	470 
    -- CP-element group 472: successors 
    -- CP-element group 472: marked-successors 
    -- CP-element group 472: 	443 
    -- CP-element group 472: 	451 
    -- CP-element group 472: 	470 
    -- CP-element group 472:  members (3) 
      -- CP-element group 472: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_965_sample_completed_
      -- CP-element group 472: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_965_Sample/$exit
      -- CP-element group 472: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_965_Sample/ack
      -- 
    ack_2065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 472_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue219_exec_guard_894_delayed_1_0_963_inst_ack_0, ack => zeropad_CP_182_elements(472)); -- 
    -- CP-element group 473:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	471 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	611 
    -- CP-element group 473: marked-successors 
    -- CP-element group 473: 	471 
    -- CP-element group 473:  members (3) 
      -- CP-element group 473: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_965_update_completed_
      -- CP-element group 473: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_965_Update/$exit
      -- CP-element group 473: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_965_Update/ack
      -- 
    ack_2070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 473_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue219_exec_guard_894_delayed_1_0_963_inst_ack_1, ack => zeropad_CP_182_elements(473)); -- 
    -- CP-element group 474:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	445 
    -- CP-element group 474: 	453 
    -- CP-element group 474: marked-predecessors 
    -- CP-element group 474: 	476 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	476 
    -- CP-element group 474:  members (3) 
      -- CP-element group 474: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_974_sample_start_
      -- CP-element group 474: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_974_Sample/$entry
      -- CP-element group 474: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_974_Sample/req
      -- 
    req_2078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(474), ack => W_landx_xlhsx_xtrue219_exec_guard_900_delayed_1_0_972_inst_req_0); -- 
    zeropad_cp_element_group_474: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_474"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(445) & zeropad_CP_182_elements(453) & zeropad_CP_182_elements(476);
      gj_zeropad_cp_element_group_474 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(474), clk => clk, reset => reset); --
    end block;
    -- CP-element group 475:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: marked-predecessors 
    -- CP-element group 475: 	477 
    -- CP-element group 475: successors 
    -- CP-element group 475: 	477 
    -- CP-element group 475:  members (3) 
      -- CP-element group 475: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_974_update_start_
      -- CP-element group 475: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_974_Update/$entry
      -- CP-element group 475: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_974_Update/req
      -- 
    req_2083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(475), ack => W_landx_xlhsx_xtrue219_exec_guard_900_delayed_1_0_972_inst_req_1); -- 
    zeropad_cp_element_group_475: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_475"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_CP_182_elements(477);
      gj_zeropad_cp_element_group_475 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(475), clk => clk, reset => reset); --
    end block;
    -- CP-element group 476:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	474 
    -- CP-element group 476: successors 
    -- CP-element group 476: marked-successors 
    -- CP-element group 476: 	443 
    -- CP-element group 476: 	451 
    -- CP-element group 476: 	474 
    -- CP-element group 476:  members (3) 
      -- CP-element group 476: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_974_sample_completed_
      -- CP-element group 476: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_974_Sample/$exit
      -- CP-element group 476: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_974_Sample/ack
      -- 
    ack_2079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 476_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue219_exec_guard_900_delayed_1_0_972_inst_ack_0, ack => zeropad_CP_182_elements(476)); -- 
    -- CP-element group 477:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	475 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	611 
    -- CP-element group 477: marked-successors 
    -- CP-element group 477: 	475 
    -- CP-element group 477:  members (3) 
      -- CP-element group 477: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_974_update_completed_
      -- CP-element group 477: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_974_Update/$exit
      -- CP-element group 477: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_974_Update/ack
      -- 
    ack_2084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 477_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue219_exec_guard_900_delayed_1_0_972_inst_ack_1, ack => zeropad_CP_182_elements(477)); -- 
    -- CP-element group 478:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	469 
    -- CP-element group 478: marked-predecessors 
    -- CP-element group 478: 	480 
    -- CP-element group 478: successors 
    -- CP-element group 478: 	480 
    -- CP-element group 478:  members (3) 
      -- CP-element group 478: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_977_sample_start_
      -- CP-element group 478: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_977_Sample/$entry
      -- CP-element group 478: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_977_Sample/req
      -- 
    req_2092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(478), ack => W_add234_903_delayed_1_0_975_inst_req_0); -- 
    zeropad_cp_element_group_478: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_478"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(469) & zeropad_CP_182_elements(480);
      gj_zeropad_cp_element_group_478 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(478), clk => clk, reset => reset); --
    end block;
    -- CP-element group 479:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	115 
    -- CP-element group 479: marked-predecessors 
    -- CP-element group 479: 	481 
    -- CP-element group 479: successors 
    -- CP-element group 479: 	481 
    -- CP-element group 479:  members (3) 
      -- CP-element group 479: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_977_update_start_
      -- CP-element group 479: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_977_Update/$entry
      -- CP-element group 479: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_977_Update/req
      -- 
    req_2097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(479), ack => W_add234_903_delayed_1_0_975_inst_req_1); -- 
    zeropad_cp_element_group_479: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_479"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(481);
      gj_zeropad_cp_element_group_479 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(479), clk => clk, reset => reset); --
    end block;
    -- CP-element group 480:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	478 
    -- CP-element group 480: successors 
    -- CP-element group 480: marked-successors 
    -- CP-element group 480: 	467 
    -- CP-element group 480: 	478 
    -- CP-element group 480:  members (3) 
      -- CP-element group 480: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_977_sample_completed_
      -- CP-element group 480: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_977_Sample/$exit
      -- CP-element group 480: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_977_Sample/ack
      -- 
    ack_2093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 480_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add234_903_delayed_1_0_975_inst_ack_0, ack => zeropad_CP_182_elements(480)); -- 
    -- CP-element group 481:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	479 
    -- CP-element group 481: successors 
    -- CP-element group 481: 	611 
    -- CP-element group 481: marked-successors 
    -- CP-element group 481: 	137 
    -- CP-element group 481: 	479 
    -- CP-element group 481:  members (3) 
      -- CP-element group 481: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_977_update_completed_
      -- CP-element group 481: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_977_Update/$exit
      -- CP-element group 481: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_977_Update/ack
      -- 
    ack_2098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 481_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add234_903_delayed_1_0_975_inst_ack_1, ack => zeropad_CP_182_elements(481)); -- 
    -- CP-element group 482:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	142 
    -- CP-element group 482: marked-predecessors 
    -- CP-element group 482: 	484 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	484 
    -- CP-element group 482:  members (3) 
      -- CP-element group 482: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_980_sample_start_
      -- CP-element group 482: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_980_Sample/$entry
      -- CP-element group 482: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_980_Sample/req
      -- 
    req_2106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(482), ack => W_target_out_offsetx_x1_904_delayed_3_0_978_inst_req_0); -- 
    zeropad_cp_element_group_482: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_482"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(484);
      gj_zeropad_cp_element_group_482 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(482), clk => clk, reset => reset); --
    end block;
    -- CP-element group 483:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	115 
    -- CP-element group 483: marked-predecessors 
    -- CP-element group 483: 	485 
    -- CP-element group 483: successors 
    -- CP-element group 483: 	485 
    -- CP-element group 483:  members (3) 
      -- CP-element group 483: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_980_update_start_
      -- CP-element group 483: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_980_Update/$entry
      -- CP-element group 483: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_980_Update/req
      -- 
    req_2111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(483), ack => W_target_out_offsetx_x1_904_delayed_3_0_978_inst_req_1); -- 
    zeropad_cp_element_group_483: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_483"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(485);
      gj_zeropad_cp_element_group_483 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(483), clk => clk, reset => reset); --
    end block;
    -- CP-element group 484:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	482 
    -- CP-element group 484: successors 
    -- CP-element group 484: marked-successors 
    -- CP-element group 484: 	138 
    -- CP-element group 484: 	482 
    -- CP-element group 484:  members (3) 
      -- CP-element group 484: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_980_sample_completed_
      -- CP-element group 484: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_980_Sample/$exit
      -- CP-element group 484: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_980_Sample/ack
      -- 
    ack_2107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 484_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_target_out_offsetx_x1_904_delayed_3_0_978_inst_ack_0, ack => zeropad_CP_182_elements(484)); -- 
    -- CP-element group 485:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	483 
    -- CP-element group 485: successors 
    -- CP-element group 485: 	611 
    -- CP-element group 485: marked-successors 
    -- CP-element group 485: 	137 
    -- CP-element group 485: 	483 
    -- CP-element group 485:  members (3) 
      -- CP-element group 485: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_980_update_completed_
      -- CP-element group 485: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_980_Update/$exit
      -- CP-element group 485: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_980_Update/ack
      -- 
    ack_2112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 485_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_target_out_offsetx_x1_904_delayed_3_0_978_inst_ack_1, ack => zeropad_CP_182_elements(485)); -- 
    -- CP-element group 486:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: 	413 
    -- CP-element group 486: 	425 
    -- CP-element group 486: 	433 
    -- CP-element group 486: marked-predecessors 
    -- CP-element group 486: 	488 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	488 
    -- CP-element group 486:  members (3) 
      -- CP-element group 486: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_993_sample_start_
      -- CP-element group 486: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_993_Sample/$entry
      -- CP-element group 486: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_993_Sample/req
      -- 
    req_2120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(486), ack => W_ifx_xthen191_condx_xend_taken_911_delayed_1_0_991_inst_req_0); -- 
    zeropad_cp_element_group_486: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_486"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(413) & zeropad_CP_182_elements(425) & zeropad_CP_182_elements(433) & zeropad_CP_182_elements(488);
      gj_zeropad_cp_element_group_486 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(486), clk => clk, reset => reset); --
    end block;
    -- CP-element group 487:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	115 
    -- CP-element group 487: marked-predecessors 
    -- CP-element group 487: 	489 
    -- CP-element group 487: 	512 
    -- CP-element group 487: 	520 
    -- CP-element group 487: 	548 
    -- CP-element group 487: 	571 
    -- CP-element group 487: successors 
    -- CP-element group 487: 	489 
    -- CP-element group 487:  members (3) 
      -- CP-element group 487: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_993_update_start_
      -- CP-element group 487: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_993_Update/$entry
      -- CP-element group 487: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_993_Update/req
      -- 
    req_2125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(487), ack => W_ifx_xthen191_condx_xend_taken_911_delayed_1_0_991_inst_req_1); -- 
    zeropad_cp_element_group_487: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_487"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(489) & zeropad_CP_182_elements(512) & zeropad_CP_182_elements(520) & zeropad_CP_182_elements(548) & zeropad_CP_182_elements(571);
      gj_zeropad_cp_element_group_487 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(487), clk => clk, reset => reset); --
    end block;
    -- CP-element group 488:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	486 
    -- CP-element group 488: successors 
    -- CP-element group 488: marked-successors 
    -- CP-element group 488: 	411 
    -- CP-element group 488: 	423 
    -- CP-element group 488: 	431 
    -- CP-element group 488: 	486 
    -- CP-element group 488:  members (3) 
      -- CP-element group 488: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_993_sample_completed_
      -- CP-element group 488: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_993_Sample/$exit
      -- CP-element group 488: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_993_Sample/ack
      -- 
    ack_2121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 488_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen191_condx_xend_taken_911_delayed_1_0_991_inst_ack_0, ack => zeropad_CP_182_elements(488)); -- 
    -- CP-element group 489:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	487 
    -- CP-element group 489: successors 
    -- CP-element group 489: 	510 
    -- CP-element group 489: 	518 
    -- CP-element group 489: 	546 
    -- CP-element group 489: 	569 
    -- CP-element group 489: marked-successors 
    -- CP-element group 489: 	118 
    -- CP-element group 489: 	179 
    -- CP-element group 489: 	200 
    -- CP-element group 489: 	221 
    -- CP-element group 489: 	305 
    -- CP-element group 489: 	487 
    -- CP-element group 489:  members (3) 
      -- CP-element group 489: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_993_update_completed_
      -- CP-element group 489: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_993_Update/$exit
      -- CP-element group 489: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_993_Update/ack
      -- 
    ack_2126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 489_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen191_condx_xend_taken_911_delayed_1_0_991_inst_ack_1, ack => zeropad_CP_182_elements(489)); -- 
    -- CP-element group 490:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: 	413 
    -- CP-element group 490: 	425 
    -- CP-element group 490: 	433 
    -- CP-element group 490: marked-predecessors 
    -- CP-element group 490: 	492 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	492 
    -- CP-element group 490:  members (3) 
      -- CP-element group 490: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1003_sample_start_
      -- CP-element group 490: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1003_Sample/$entry
      -- CP-element group 490: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1003_Sample/req
      -- 
    req_2134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(490), ack => W_ifx_xthen191_condx_xend_taken_918_delayed_2_0_1001_inst_req_0); -- 
    zeropad_cp_element_group_490: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_490"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(413) & zeropad_CP_182_elements(425) & zeropad_CP_182_elements(433) & zeropad_CP_182_elements(492);
      gj_zeropad_cp_element_group_490 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(490), clk => clk, reset => reset); --
    end block;
    -- CP-element group 491:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	115 
    -- CP-element group 491: marked-predecessors 
    -- CP-element group 491: 	493 
    -- CP-element group 491: successors 
    -- CP-element group 491: 	493 
    -- CP-element group 491:  members (3) 
      -- CP-element group 491: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1003_update_start_
      -- CP-element group 491: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1003_Update/$entry
      -- CP-element group 491: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1003_Update/req
      -- 
    req_2139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(491), ack => W_ifx_xthen191_condx_xend_taken_918_delayed_2_0_1001_inst_req_1); -- 
    zeropad_cp_element_group_491: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_491"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(493);
      gj_zeropad_cp_element_group_491 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(491), clk => clk, reset => reset); --
    end block;
    -- CP-element group 492:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	490 
    -- CP-element group 492: successors 
    -- CP-element group 492: marked-successors 
    -- CP-element group 492: 	411 
    -- CP-element group 492: 	423 
    -- CP-element group 492: 	431 
    -- CP-element group 492: 	490 
    -- CP-element group 492:  members (3) 
      -- CP-element group 492: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1003_sample_completed_
      -- CP-element group 492: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1003_Sample/$exit
      -- CP-element group 492: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1003_Sample/ack
      -- 
    ack_2135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen191_condx_xend_taken_918_delayed_2_0_1001_inst_ack_0, ack => zeropad_CP_182_elements(492)); -- 
    -- CP-element group 493:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	491 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	611 
    -- CP-element group 493: marked-successors 
    -- CP-element group 493: 	137 
    -- CP-element group 493: 	491 
    -- CP-element group 493:  members (3) 
      -- CP-element group 493: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1003_update_completed_
      -- CP-element group 493: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1003_Update/$exit
      -- CP-element group 493: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1003_Update/ack
      -- 
    ack_2140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 493_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen191_condx_xend_taken_918_delayed_2_0_1001_inst_ack_1, ack => zeropad_CP_182_elements(493)); -- 
    -- CP-element group 494:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	142 
    -- CP-element group 494: marked-predecessors 
    -- CP-element group 494: 	496 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	496 
    -- CP-element group 494:  members (3) 
      -- CP-element group 494: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1006_sample_start_
      -- CP-element group 494: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1006_Sample/$entry
      -- CP-element group 494: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1006_Sample/rr
      -- 
    rr_2148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(494), ack => type_cast_1006_inst_req_0); -- 
    zeropad_cp_element_group_494: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_494"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(496);
      gj_zeropad_cp_element_group_494 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(494), clk => clk, reset => reset); --
    end block;
    -- CP-element group 495:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	115 
    -- CP-element group 495: marked-predecessors 
    -- CP-element group 495: 	497 
    -- CP-element group 495: successors 
    -- CP-element group 495: 	497 
    -- CP-element group 495:  members (3) 
      -- CP-element group 495: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1006_update_start_
      -- CP-element group 495: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1006_Update/$entry
      -- CP-element group 495: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1006_Update/cr
      -- 
    cr_2153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(495), ack => type_cast_1006_inst_req_1); -- 
    zeropad_cp_element_group_495: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_495"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(497);
      gj_zeropad_cp_element_group_495 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(495), clk => clk, reset => reset); --
    end block;
    -- CP-element group 496:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	494 
    -- CP-element group 496: successors 
    -- CP-element group 496: marked-successors 
    -- CP-element group 496: 	138 
    -- CP-element group 496: 	494 
    -- CP-element group 496:  members (3) 
      -- CP-element group 496: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1006_sample_completed_
      -- CP-element group 496: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1006_Sample/$exit
      -- CP-element group 496: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1006_Sample/ra
      -- 
    ra_2149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 496_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1006_inst_ack_0, ack => zeropad_CP_182_elements(496)); -- 
    -- CP-element group 497:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: 	495 
    -- CP-element group 497: successors 
    -- CP-element group 497: 	611 
    -- CP-element group 497: marked-successors 
    -- CP-element group 497: 	137 
    -- CP-element group 497: 	495 
    -- CP-element group 497:  members (3) 
      -- CP-element group 497: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1006_update_completed_
      -- CP-element group 497: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1006_Update/$exit
      -- CP-element group 497: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1006_Update/ca
      -- 
    ca_2154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 497_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1006_inst_ack_1, ack => zeropad_CP_182_elements(497)); -- 
    -- CP-element group 498:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 498: predecessors 
    -- CP-element group 498: 	445 
    -- CP-element group 498: 	457 
    -- CP-element group 498: marked-predecessors 
    -- CP-element group 498: 	500 
    -- CP-element group 498: successors 
    -- CP-element group 498: 	500 
    -- CP-element group 498:  members (3) 
      -- CP-element group 498: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1010_sample_start_
      -- CP-element group 498: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1010_Sample/$entry
      -- CP-element group 498: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1010_Sample/req
      -- 
    req_2162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(498), ack => W_landx_xlhsx_xtrue208_condx_xend_taken_921_delayed_1_0_1008_inst_req_0); -- 
    zeropad_cp_element_group_498: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_498"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(445) & zeropad_CP_182_elements(457) & zeropad_CP_182_elements(500);
      gj_zeropad_cp_element_group_498 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(498), clk => clk, reset => reset); --
    end block;
    -- CP-element group 499:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 499: predecessors 
    -- CP-element group 499: 	115 
    -- CP-element group 499: marked-predecessors 
    -- CP-element group 499: 	501 
    -- CP-element group 499: successors 
    -- CP-element group 499: 	501 
    -- CP-element group 499:  members (3) 
      -- CP-element group 499: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1010_update_start_
      -- CP-element group 499: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1010_Update/$entry
      -- CP-element group 499: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1010_Update/req
      -- 
    req_2167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(499), ack => W_landx_xlhsx_xtrue208_condx_xend_taken_921_delayed_1_0_1008_inst_req_1); -- 
    zeropad_cp_element_group_499: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_499"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(501);
      gj_zeropad_cp_element_group_499 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(499), clk => clk, reset => reset); --
    end block;
    -- CP-element group 500:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 500: predecessors 
    -- CP-element group 500: 	498 
    -- CP-element group 500: successors 
    -- CP-element group 500: marked-successors 
    -- CP-element group 500: 	443 
    -- CP-element group 500: 	455 
    -- CP-element group 500: 	498 
    -- CP-element group 500:  members (3) 
      -- CP-element group 500: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1010_sample_completed_
      -- CP-element group 500: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1010_Sample/$exit
      -- CP-element group 500: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1010_Sample/ack
      -- 
    ack_2163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 500_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue208_condx_xend_taken_921_delayed_1_0_1008_inst_ack_0, ack => zeropad_CP_182_elements(500)); -- 
    -- CP-element group 501:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 501: predecessors 
    -- CP-element group 501: 	499 
    -- CP-element group 501: successors 
    -- CP-element group 501: 	611 
    -- CP-element group 501: marked-successors 
    -- CP-element group 501: 	137 
    -- CP-element group 501: 	499 
    -- CP-element group 501:  members (3) 
      -- CP-element group 501: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1010_update_completed_
      -- CP-element group 501: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1010_Update/$exit
      -- CP-element group 501: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1010_Update/ack
      -- 
    ack_2168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 501_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue208_condx_xend_taken_921_delayed_1_0_1008_inst_ack_1, ack => zeropad_CP_182_elements(501)); -- 
    -- CP-element group 502:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 502: predecessors 
    -- CP-element group 502: 	142 
    -- CP-element group 502: marked-predecessors 
    -- CP-element group 502: 	504 
    -- CP-element group 502: successors 
    -- CP-element group 502: 	504 
    -- CP-element group 502:  members (3) 
      -- CP-element group 502: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1013_sample_start_
      -- CP-element group 502: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1013_Sample/$entry
      -- CP-element group 502: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1013_Sample/rr
      -- 
    rr_2176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(502), ack => type_cast_1013_inst_req_0); -- 
    zeropad_cp_element_group_502: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_502"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(504);
      gj_zeropad_cp_element_group_502 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(502), clk => clk, reset => reset); --
    end block;
    -- CP-element group 503:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 503: predecessors 
    -- CP-element group 503: 	115 
    -- CP-element group 503: marked-predecessors 
    -- CP-element group 503: 	505 
    -- CP-element group 503: successors 
    -- CP-element group 503: 	505 
    -- CP-element group 503:  members (3) 
      -- CP-element group 503: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1013_update_start_
      -- CP-element group 503: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1013_Update/$entry
      -- CP-element group 503: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1013_Update/cr
      -- 
    cr_2181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(503), ack => type_cast_1013_inst_req_1); -- 
    zeropad_cp_element_group_503: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_503"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(505);
      gj_zeropad_cp_element_group_503 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(503), clk => clk, reset => reset); --
    end block;
    -- CP-element group 504:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 504: predecessors 
    -- CP-element group 504: 	502 
    -- CP-element group 504: successors 
    -- CP-element group 504: marked-successors 
    -- CP-element group 504: 	138 
    -- CP-element group 504: 	502 
    -- CP-element group 504:  members (3) 
      -- CP-element group 504: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1013_sample_completed_
      -- CP-element group 504: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1013_Sample/$exit
      -- CP-element group 504: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1013_Sample/ra
      -- 
    ra_2177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 504_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1013_inst_ack_0, ack => zeropad_CP_182_elements(504)); -- 
    -- CP-element group 505:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 505: predecessors 
    -- CP-element group 505: 	503 
    -- CP-element group 505: successors 
    -- CP-element group 505: 	611 
    -- CP-element group 505: marked-successors 
    -- CP-element group 505: 	137 
    -- CP-element group 505: 	503 
    -- CP-element group 505:  members (3) 
      -- CP-element group 505: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1013_update_completed_
      -- CP-element group 505: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1013_Update/$exit
      -- CP-element group 505: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1013_Update/ca
      -- 
    ca_2182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 505_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1013_inst_ack_1, ack => zeropad_CP_182_elements(505)); -- 
    -- CP-element group 506:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 506: predecessors 
    -- CP-element group 506: 	445 
    -- CP-element group 506: 	453 
    -- CP-element group 506: marked-predecessors 
    -- CP-element group 506: 	508 
    -- CP-element group 506: successors 
    -- CP-element group 506: 	508 
    -- CP-element group 506:  members (3) 
      -- CP-element group 506: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1017_sample_start_
      -- CP-element group 506: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1017_Sample/$entry
      -- CP-element group 506: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1017_Sample/req
      -- 
    req_2190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(506), ack => W_landx_xlhsx_xtrue219_condx_xend_taken_924_delayed_1_0_1015_inst_req_0); -- 
    zeropad_cp_element_group_506: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_506"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(445) & zeropad_CP_182_elements(453) & zeropad_CP_182_elements(508);
      gj_zeropad_cp_element_group_506 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(506), clk => clk, reset => reset); --
    end block;
    -- CP-element group 507:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 507: predecessors 
    -- CP-element group 507: 	115 
    -- CP-element group 507: marked-predecessors 
    -- CP-element group 507: 	509 
    -- CP-element group 507: successors 
    -- CP-element group 507: 	509 
    -- CP-element group 507:  members (3) 
      -- CP-element group 507: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1017_update_start_
      -- CP-element group 507: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1017_Update/$entry
      -- CP-element group 507: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1017_Update/req
      -- 
    req_2195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(507), ack => W_landx_xlhsx_xtrue219_condx_xend_taken_924_delayed_1_0_1015_inst_req_1); -- 
    zeropad_cp_element_group_507: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_507"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(509);
      gj_zeropad_cp_element_group_507 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(507), clk => clk, reset => reset); --
    end block;
    -- CP-element group 508:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 508: predecessors 
    -- CP-element group 508: 	506 
    -- CP-element group 508: successors 
    -- CP-element group 508: marked-successors 
    -- CP-element group 508: 	443 
    -- CP-element group 508: 	451 
    -- CP-element group 508: 	506 
    -- CP-element group 508:  members (3) 
      -- CP-element group 508: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1017_sample_completed_
      -- CP-element group 508: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1017_Sample/$exit
      -- CP-element group 508: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1017_Sample/ack
      -- 
    ack_2191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 508_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue219_condx_xend_taken_924_delayed_1_0_1015_inst_ack_0, ack => zeropad_CP_182_elements(508)); -- 
    -- CP-element group 509:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 509: predecessors 
    -- CP-element group 509: 	507 
    -- CP-element group 509: successors 
    -- CP-element group 509: 	611 
    -- CP-element group 509: marked-successors 
    -- CP-element group 509: 	137 
    -- CP-element group 509: 	507 
    -- CP-element group 509:  members (3) 
      -- CP-element group 509: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1017_update_completed_
      -- CP-element group 509: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1017_Update/$exit
      -- CP-element group 509: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1017_Update/ack
      -- 
    ack_2196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 509_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_landx_xlhsx_xtrue219_condx_xend_taken_924_delayed_1_0_1015_inst_ack_1, ack => zeropad_CP_182_elements(509)); -- 
    -- CP-element group 510:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 510: predecessors 
    -- CP-element group 510: 	445 
    -- CP-element group 510: 	453 
    -- CP-element group 510: 	457 
    -- CP-element group 510: 	489 
    -- CP-element group 510: marked-predecessors 
    -- CP-element group 510: 	512 
    -- CP-element group 510: successors 
    -- CP-element group 510: 	512 
    -- CP-element group 510:  members (3) 
      -- CP-element group 510: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1034_sample_start_
      -- CP-element group 510: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1034_Sample/$entry
      -- CP-element group 510: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1034_Sample/req
      -- 
    req_2204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(510), ack => W_condx_xend_exec_guard_933_delayed_1_0_1032_inst_req_0); -- 
    zeropad_cp_element_group_510: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_510"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(445) & zeropad_CP_182_elements(453) & zeropad_CP_182_elements(457) & zeropad_CP_182_elements(489) & zeropad_CP_182_elements(512);
      gj_zeropad_cp_element_group_510 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(510), clk => clk, reset => reset); --
    end block;
    -- CP-element group 511:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 511: predecessors 
    -- CP-element group 511: marked-predecessors 
    -- CP-element group 511: 	513 
    -- CP-element group 511: successors 
    -- CP-element group 511: 	513 
    -- CP-element group 511:  members (3) 
      -- CP-element group 511: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1034_update_start_
      -- CP-element group 511: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1034_Update/$entry
      -- CP-element group 511: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1034_Update/req
      -- 
    req_2209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(511), ack => W_condx_xend_exec_guard_933_delayed_1_0_1032_inst_req_1); -- 
    zeropad_cp_element_group_511: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_511"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_CP_182_elements(513);
      gj_zeropad_cp_element_group_511 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(511), clk => clk, reset => reset); --
    end block;
    -- CP-element group 512:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 512: predecessors 
    -- CP-element group 512: 	510 
    -- CP-element group 512: successors 
    -- CP-element group 512: marked-successors 
    -- CP-element group 512: 	443 
    -- CP-element group 512: 	451 
    -- CP-element group 512: 	455 
    -- CP-element group 512: 	487 
    -- CP-element group 512: 	510 
    -- CP-element group 512:  members (3) 
      -- CP-element group 512: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1034_sample_completed_
      -- CP-element group 512: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1034_Sample/$exit
      -- CP-element group 512: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1034_Sample/ack
      -- 
    ack_2205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 512_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_condx_xend_exec_guard_933_delayed_1_0_1032_inst_ack_0, ack => zeropad_CP_182_elements(512)); -- 
    -- CP-element group 513:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 513: predecessors 
    -- CP-element group 513: 	511 
    -- CP-element group 513: successors 
    -- CP-element group 513: 	611 
    -- CP-element group 513: marked-successors 
    -- CP-element group 513: 	511 
    -- CP-element group 513:  members (3) 
      -- CP-element group 513: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1034_update_completed_
      -- CP-element group 513: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1034_Update/$exit
      -- CP-element group 513: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1034_Update/ack
      -- 
    ack_2210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 513_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_condx_xend_exec_guard_933_delayed_1_0_1032_inst_ack_1, ack => zeropad_CP_182_elements(513)); -- 
    -- CP-element group 514:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 514: predecessors 
    -- CP-element group 514: 	142 
    -- CP-element group 514: 	163 
    -- CP-element group 514: marked-predecessors 
    -- CP-element group 514: 	516 
    -- CP-element group 514: successors 
    -- CP-element group 514: 	516 
    -- CP-element group 514:  members (3) 
      -- CP-element group 514: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1047_sample_start_
      -- CP-element group 514: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1047_Sample/$entry
      -- CP-element group 514: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1047_Sample/req
      -- 
    req_2218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(514), ack => W_ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1045_inst_req_0); -- 
    zeropad_cp_element_group_514: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_514"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(516);
      gj_zeropad_cp_element_group_514 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(514), clk => clk, reset => reset); --
    end block;
    -- CP-element group 515:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 515: predecessors 
    -- CP-element group 515: 	115 
    -- CP-element group 515: marked-predecessors 
    -- CP-element group 515: 	517 
    -- CP-element group 515: successors 
    -- CP-element group 515: 	517 
    -- CP-element group 515:  members (3) 
      -- CP-element group 515: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1047_update_start_
      -- CP-element group 515: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1047_Update/$entry
      -- CP-element group 515: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1047_Update/req
      -- 
    req_2223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(515), ack => W_ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1045_inst_req_1); -- 
    zeropad_cp_element_group_515: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_515"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(517);
      gj_zeropad_cp_element_group_515 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(515), clk => clk, reset => reset); --
    end block;
    -- CP-element group 516:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 516: predecessors 
    -- CP-element group 516: 	514 
    -- CP-element group 516: successors 
    -- CP-element group 516: marked-successors 
    -- CP-element group 516: 	138 
    -- CP-element group 516: 	159 
    -- CP-element group 516: 	514 
    -- CP-element group 516:  members (3) 
      -- CP-element group 516: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1047_sample_completed_
      -- CP-element group 516: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1047_Sample/$exit
      -- CP-element group 516: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1047_Sample/ack
      -- 
    ack_2219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 516_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1045_inst_ack_0, ack => zeropad_CP_182_elements(516)); -- 
    -- CP-element group 517:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 517: predecessors 
    -- CP-element group 517: 	515 
    -- CP-element group 517: successors 
    -- CP-element group 517: 	611 
    -- CP-element group 517: marked-successors 
    -- CP-element group 517: 	179 
    -- CP-element group 517: 	200 
    -- CP-element group 517: 	305 
    -- CP-element group 517: 	515 
    -- CP-element group 517:  members (3) 
      -- CP-element group 517: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1047_update_completed_
      -- CP-element group 517: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1047_Update/$exit
      -- CP-element group 517: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1047_Update/ack
      -- 
    ack_2224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 517_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1045_inst_ack_1, ack => zeropad_CP_182_elements(517)); -- 
    -- CP-element group 518:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 518: predecessors 
    -- CP-element group 518: 	445 
    -- CP-element group 518: 	453 
    -- CP-element group 518: 	457 
    -- CP-element group 518: 	489 
    -- CP-element group 518: marked-predecessors 
    -- CP-element group 518: 	520 
    -- CP-element group 518: successors 
    -- CP-element group 518: 	520 
    -- CP-element group 518:  members (3) 
      -- CP-element group 518: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1055_sample_start_
      -- CP-element group 518: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1055_Sample/$entry
      -- CP-element group 518: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1055_Sample/req
      -- 
    req_2232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(518), ack => W_condx_xend_ifx_xend238_taken_949_delayed_10_0_1053_inst_req_0); -- 
    zeropad_cp_element_group_518: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_518"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(445) & zeropad_CP_182_elements(453) & zeropad_CP_182_elements(457) & zeropad_CP_182_elements(489) & zeropad_CP_182_elements(520);
      gj_zeropad_cp_element_group_518 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(518), clk => clk, reset => reset); --
    end block;
    -- CP-element group 519:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 519: predecessors 
    -- CP-element group 519: 	115 
    -- CP-element group 519: marked-predecessors 
    -- CP-element group 519: 	521 
    -- CP-element group 519: successors 
    -- CP-element group 519: 	521 
    -- CP-element group 519:  members (3) 
      -- CP-element group 519: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1055_update_start_
      -- CP-element group 519: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1055_Update/$entry
      -- CP-element group 519: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1055_Update/req
      -- 
    req_2237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(519), ack => W_condx_xend_ifx_xend238_taken_949_delayed_10_0_1053_inst_req_1); -- 
    zeropad_cp_element_group_519: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_519"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(521);
      gj_zeropad_cp_element_group_519 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(519), clk => clk, reset => reset); --
    end block;
    -- CP-element group 520:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 520: predecessors 
    -- CP-element group 520: 	518 
    -- CP-element group 520: successors 
    -- CP-element group 520: marked-successors 
    -- CP-element group 520: 	443 
    -- CP-element group 520: 	451 
    -- CP-element group 520: 	455 
    -- CP-element group 520: 	487 
    -- CP-element group 520: 	518 
    -- CP-element group 520:  members (3) 
      -- CP-element group 520: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1055_sample_completed_
      -- CP-element group 520: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1055_Sample/$exit
      -- CP-element group 520: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1055_Sample/ack
      -- 
    ack_2233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 520_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_condx_xend_ifx_xend238_taken_949_delayed_10_0_1053_inst_ack_0, ack => zeropad_CP_182_elements(520)); -- 
    -- CP-element group 521:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 521: predecessors 
    -- CP-element group 521: 	519 
    -- CP-element group 521: successors 
    -- CP-element group 521: 	611 
    -- CP-element group 521: marked-successors 
    -- CP-element group 521: 	326 
    -- CP-element group 521: 	519 
    -- CP-element group 521:  members (3) 
      -- CP-element group 521: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1055_update_completed_
      -- CP-element group 521: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1055_Update/$exit
      -- CP-element group 521: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1055_Update/ack
      -- 
    ack_2238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 521_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_condx_xend_ifx_xend238_taken_949_delayed_10_0_1053_inst_ack_1, ack => zeropad_CP_182_elements(521)); -- 
    -- CP-element group 522:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 522: predecessors 
    -- CP-element group 522: 	142 
    -- CP-element group 522: 	163 
    -- CP-element group 522: 	331 
    -- CP-element group 522: marked-predecessors 
    -- CP-element group 522: 	524 
    -- CP-element group 522: successors 
    -- CP-element group 522: 	524 
    -- CP-element group 522:  members (3) 
      -- CP-element group 522: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1062_sample_start_
      -- CP-element group 522: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1062_start/$entry
      -- CP-element group 522: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1062_start/req
      -- 
    req_2246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(522), ack => MUX_1062_inst_req_0); -- 
    zeropad_cp_element_group_522: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_522"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(331) & zeropad_CP_182_elements(524);
      gj_zeropad_cp_element_group_522 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(522), clk => clk, reset => reset); --
    end block;
    -- CP-element group 523:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 523: predecessors 
    -- CP-element group 523: 	115 
    -- CP-element group 523: marked-predecessors 
    -- CP-element group 523: 	525 
    -- CP-element group 523: successors 
    -- CP-element group 523: 	525 
    -- CP-element group 523:  members (3) 
      -- CP-element group 523: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1062_update_start_
      -- CP-element group 523: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1062_complete/$entry
      -- CP-element group 523: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1062_complete/req
      -- 
    req_2251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(523), ack => MUX_1062_inst_req_1); -- 
    zeropad_cp_element_group_523: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_523"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(525);
      gj_zeropad_cp_element_group_523 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(523), clk => clk, reset => reset); --
    end block;
    -- CP-element group 524:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 524: predecessors 
    -- CP-element group 524: 	522 
    -- CP-element group 524: successors 
    -- CP-element group 524: marked-successors 
    -- CP-element group 524: 	138 
    -- CP-element group 524: 	159 
    -- CP-element group 524: 	327 
    -- CP-element group 524: 	522 
    -- CP-element group 524:  members (3) 
      -- CP-element group 524: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1062_sample_completed_
      -- CP-element group 524: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1062_start/$exit
      -- CP-element group 524: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1062_start/ack
      -- 
    ack_2247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 524_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1062_inst_ack_0, ack => zeropad_CP_182_elements(524)); -- 
    -- CP-element group 525:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 525: predecessors 
    -- CP-element group 525: 	523 
    -- CP-element group 525: successors 
    -- CP-element group 525: 	611 
    -- CP-element group 525: marked-successors 
    -- CP-element group 525: 	326 
    -- CP-element group 525: 	523 
    -- CP-element group 525:  members (3) 
      -- CP-element group 525: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1062_update_completed_
      -- CP-element group 525: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1062_complete/$exit
      -- CP-element group 525: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1062_complete/ack
      -- 
    ack_2252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 525_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1062_inst_ack_1, ack => zeropad_CP_182_elements(525)); -- 
    -- CP-element group 526:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 526: predecessors 
    -- CP-element group 526: 	142 
    -- CP-element group 526: 	163 
    -- CP-element group 526: 	226 
    -- CP-element group 526: marked-predecessors 
    -- CP-element group 526: 	528 
    -- CP-element group 526: successors 
    -- CP-element group 526: 	528 
    -- CP-element group 526:  members (3) 
      -- CP-element group 526: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1073_sample_start_
      -- CP-element group 526: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1073_Sample/$entry
      -- CP-element group 526: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1073_Sample/rr
      -- 
    rr_2260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(526), ack => type_cast_1073_inst_req_0); -- 
    zeropad_cp_element_group_526: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_526"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(226) & zeropad_CP_182_elements(528);
      gj_zeropad_cp_element_group_526 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(526), clk => clk, reset => reset); --
    end block;
    -- CP-element group 527:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 527: predecessors 
    -- CP-element group 527: 	115 
    -- CP-element group 527: marked-predecessors 
    -- CP-element group 527: 	529 
    -- CP-element group 527: successors 
    -- CP-element group 527: 	529 
    -- CP-element group 527:  members (3) 
      -- CP-element group 527: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1073_update_start_
      -- CP-element group 527: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1073_Update/$entry
      -- CP-element group 527: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1073_Update/cr
      -- 
    cr_2265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(527), ack => type_cast_1073_inst_req_1); -- 
    zeropad_cp_element_group_527: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_527"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(529);
      gj_zeropad_cp_element_group_527 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(527), clk => clk, reset => reset); --
    end block;
    -- CP-element group 528:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 528: predecessors 
    -- CP-element group 528: 	526 
    -- CP-element group 528: successors 
    -- CP-element group 528: marked-successors 
    -- CP-element group 528: 	138 
    -- CP-element group 528: 	159 
    -- CP-element group 528: 	222 
    -- CP-element group 528: 	526 
    -- CP-element group 528:  members (3) 
      -- CP-element group 528: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1073_sample_completed_
      -- CP-element group 528: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1073_Sample/$exit
      -- CP-element group 528: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1073_Sample/ra
      -- 
    ra_2261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 528_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1073_inst_ack_0, ack => zeropad_CP_182_elements(528)); -- 
    -- CP-element group 529:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 529: predecessors 
    -- CP-element group 529: 	527 
    -- CP-element group 529: successors 
    -- CP-element group 529: 	611 
    -- CP-element group 529: marked-successors 
    -- CP-element group 529: 	221 
    -- CP-element group 529: 	527 
    -- CP-element group 529:  members (3) 
      -- CP-element group 529: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1073_update_completed_
      -- CP-element group 529: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1073_Update/$exit
      -- CP-element group 529: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1073_Update/ca
      -- 
    ca_2266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 529_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1073_inst_ack_1, ack => zeropad_CP_182_elements(529)); -- 
    -- CP-element group 530:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 530: predecessors 
    -- CP-element group 530: 	142 
    -- CP-element group 530: 	163 
    -- CP-element group 530: 	226 
    -- CP-element group 530: marked-predecessors 
    -- CP-element group 530: 	532 
    -- CP-element group 530: successors 
    -- CP-element group 530: 	532 
    -- CP-element group 530:  members (3) 
      -- CP-element group 530: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1081_sample_start_
      -- CP-element group 530: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1081_start/$entry
      -- CP-element group 530: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1081_start/req
      -- 
    req_2274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(530), ack => MUX_1081_inst_req_0); -- 
    zeropad_cp_element_group_530: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_530"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(226) & zeropad_CP_182_elements(532);
      gj_zeropad_cp_element_group_530 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(530), clk => clk, reset => reset); --
    end block;
    -- CP-element group 531:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 531: predecessors 
    -- CP-element group 531: 	115 
    -- CP-element group 531: marked-predecessors 
    -- CP-element group 531: 	533 
    -- CP-element group 531: successors 
    -- CP-element group 531: 	533 
    -- CP-element group 531:  members (3) 
      -- CP-element group 531: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1081_update_start_
      -- CP-element group 531: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1081_complete/$entry
      -- CP-element group 531: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1081_complete/req
      -- 
    req_2279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(531), ack => MUX_1081_inst_req_1); -- 
    zeropad_cp_element_group_531: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_531"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(533);
      gj_zeropad_cp_element_group_531 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(531), clk => clk, reset => reset); --
    end block;
    -- CP-element group 532:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 532: predecessors 
    -- CP-element group 532: 	530 
    -- CP-element group 532: successors 
    -- CP-element group 532: marked-successors 
    -- CP-element group 532: 	138 
    -- CP-element group 532: 	159 
    -- CP-element group 532: 	222 
    -- CP-element group 532: 	530 
    -- CP-element group 532:  members (3) 
      -- CP-element group 532: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1081_sample_completed_
      -- CP-element group 532: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1081_start/$exit
      -- CP-element group 532: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1081_start/ack
      -- 
    ack_2275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 532_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1081_inst_ack_0, ack => zeropad_CP_182_elements(532)); -- 
    -- CP-element group 533:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 533: predecessors 
    -- CP-element group 533: 	531 
    -- CP-element group 533: successors 
    -- CP-element group 533: 	611 
    -- CP-element group 533: marked-successors 
    -- CP-element group 533: 	221 
    -- CP-element group 533: 	531 
    -- CP-element group 533:  members (3) 
      -- CP-element group 533: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1081_update_completed_
      -- CP-element group 533: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1081_complete/$exit
      -- CP-element group 533: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1081_complete/ack
      -- 
    ack_2280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 533_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1081_inst_ack_1, ack => zeropad_CP_182_elements(533)); -- 
    -- CP-element group 534:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 534: predecessors 
    -- CP-element group 534: 	121 
    -- CP-element group 534: 	142 
    -- CP-element group 534: 	163 
    -- CP-element group 534: 	226 
    -- CP-element group 534: marked-predecessors 
    -- CP-element group 534: 	536 
    -- CP-element group 534: successors 
    -- CP-element group 534: 	536 
    -- CP-element group 534:  members (3) 
      -- CP-element group 534: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1091_Sample/rr
      -- CP-element group 534: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1091_Sample/$entry
      -- CP-element group 534: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1091_sample_start_
      -- 
    rr_2288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(534), ack => type_cast_1091_inst_req_0); -- 
    zeropad_cp_element_group_534: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_534"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(121) & zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(226) & zeropad_CP_182_elements(536);
      gj_zeropad_cp_element_group_534 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(534), clk => clk, reset => reset); --
    end block;
    -- CP-element group 535:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 535: predecessors 
    -- CP-element group 535: 	115 
    -- CP-element group 535: marked-predecessors 
    -- CP-element group 535: 	537 
    -- CP-element group 535: successors 
    -- CP-element group 535: 	537 
    -- CP-element group 535:  members (3) 
      -- CP-element group 535: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1091_Update/cr
      -- CP-element group 535: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1091_Update/$entry
      -- CP-element group 535: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1091_update_start_
      -- 
    cr_2293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(535), ack => type_cast_1091_inst_req_1); -- 
    zeropad_cp_element_group_535: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_535"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(537);
      gj_zeropad_cp_element_group_535 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(535), clk => clk, reset => reset); --
    end block;
    -- CP-element group 536:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 536: predecessors 
    -- CP-element group 536: 	534 
    -- CP-element group 536: successors 
    -- CP-element group 536: marked-successors 
    -- CP-element group 536: 	119 
    -- CP-element group 536: 	138 
    -- CP-element group 536: 	159 
    -- CP-element group 536: 	222 
    -- CP-element group 536: 	534 
    -- CP-element group 536:  members (3) 
      -- CP-element group 536: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1091_Sample/ra
      -- CP-element group 536: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1091_Sample/$exit
      -- CP-element group 536: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1091_sample_completed_
      -- 
    ra_2289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 536_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1091_inst_ack_0, ack => zeropad_CP_182_elements(536)); -- 
    -- CP-element group 537:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 537: predecessors 
    -- CP-element group 537: 	535 
    -- CP-element group 537: successors 
    -- CP-element group 537: 	611 
    -- CP-element group 537: marked-successors 
    -- CP-element group 537: 	118 
    -- CP-element group 537: 	535 
    -- CP-element group 537:  members (3) 
      -- CP-element group 537: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1091_Update/ca
      -- CP-element group 537: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1091_Update/$exit
      -- CP-element group 537: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1091_update_completed_
      -- 
    ca_2294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 537_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1091_inst_ack_1, ack => zeropad_CP_182_elements(537)); -- 
    -- CP-element group 538:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 538: predecessors 
    -- CP-element group 538: 	121 
    -- CP-element group 538: 	142 
    -- CP-element group 538: 	163 
    -- CP-element group 538: marked-predecessors 
    -- CP-element group 538: 	540 
    -- CP-element group 538: successors 
    -- CP-element group 538: 	540 
    -- CP-element group 538:  members (3) 
      -- CP-element group 538: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1099_sample_start_
      -- CP-element group 538: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1099_start/$entry
      -- CP-element group 538: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1099_start/req
      -- 
    req_2302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(538), ack => MUX_1099_inst_req_0); -- 
    zeropad_cp_element_group_538: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_538"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(121) & zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(540);
      gj_zeropad_cp_element_group_538 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(538), clk => clk, reset => reset); --
    end block;
    -- CP-element group 539:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 539: predecessors 
    -- CP-element group 539: 	115 
    -- CP-element group 539: marked-predecessors 
    -- CP-element group 539: 	541 
    -- CP-element group 539: successors 
    -- CP-element group 539: 	541 
    -- CP-element group 539:  members (3) 
      -- CP-element group 539: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1099_update_start_
      -- CP-element group 539: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1099_complete/$entry
      -- CP-element group 539: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1099_complete/req
      -- 
    req_2307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(539), ack => MUX_1099_inst_req_1); -- 
    zeropad_cp_element_group_539: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_539"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(541);
      gj_zeropad_cp_element_group_539 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(539), clk => clk, reset => reset); --
    end block;
    -- CP-element group 540:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 540: predecessors 
    -- CP-element group 540: 	538 
    -- CP-element group 540: successors 
    -- CP-element group 540: marked-successors 
    -- CP-element group 540: 	119 
    -- CP-element group 540: 	138 
    -- CP-element group 540: 	159 
    -- CP-element group 540: 	538 
    -- CP-element group 540:  members (3) 
      -- CP-element group 540: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1099_sample_completed_
      -- CP-element group 540: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1099_start/$exit
      -- CP-element group 540: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1099_start/ack
      -- 
    ack_2303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 540_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1099_inst_ack_0, ack => zeropad_CP_182_elements(540)); -- 
    -- CP-element group 541:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 541: predecessors 
    -- CP-element group 541: 	539 
    -- CP-element group 541: successors 
    -- CP-element group 541: 	611 
    -- CP-element group 541: marked-successors 
    -- CP-element group 541: 	118 
    -- CP-element group 541: 	539 
    -- CP-element group 541:  members (3) 
      -- CP-element group 541: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1099_update_completed_
      -- CP-element group 541: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1099_complete/$exit
      -- CP-element group 541: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1099_complete/ack
      -- 
    ack_2308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 541_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1099_inst_ack_1, ack => zeropad_CP_182_elements(541)); -- 
    -- CP-element group 542:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 542: predecessors 
    -- CP-element group 542: 	142 
    -- CP-element group 542: 	163 
    -- CP-element group 542: 	310 
    -- CP-element group 542: marked-predecessors 
    -- CP-element group 542: 	544 
    -- CP-element group 542: successors 
    -- CP-element group 542: 	544 
    -- CP-element group 542:  members (3) 
      -- CP-element group 542: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1113_start/req
      -- CP-element group 542: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1113_start/$entry
      -- CP-element group 542: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1113_sample_start_
      -- 
    req_2316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(542), ack => MUX_1113_inst_req_0); -- 
    zeropad_cp_element_group_542: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_542"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(310) & zeropad_CP_182_elements(544);
      gj_zeropad_cp_element_group_542 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(542), clk => clk, reset => reset); --
    end block;
    -- CP-element group 543:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 543: predecessors 
    -- CP-element group 543: 	115 
    -- CP-element group 543: marked-predecessors 
    -- CP-element group 543: 	545 
    -- CP-element group 543: 	571 
    -- CP-element group 543: successors 
    -- CP-element group 543: 	545 
    -- CP-element group 543:  members (3) 
      -- CP-element group 543: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1113_complete/$entry
      -- CP-element group 543: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1113_complete/req
      -- CP-element group 543: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1113_update_start_
      -- 
    req_2321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(543), ack => MUX_1113_inst_req_1); -- 
    zeropad_cp_element_group_543: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_543"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(545) & zeropad_CP_182_elements(571);
      gj_zeropad_cp_element_group_543 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(543), clk => clk, reset => reset); --
    end block;
    -- CP-element group 544:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 544: predecessors 
    -- CP-element group 544: 	542 
    -- CP-element group 544: successors 
    -- CP-element group 544: marked-successors 
    -- CP-element group 544: 	138 
    -- CP-element group 544: 	159 
    -- CP-element group 544: 	306 
    -- CP-element group 544: 	542 
    -- CP-element group 544:  members (3) 
      -- CP-element group 544: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1113_start/$exit
      -- CP-element group 544: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1113_start/ack
      -- CP-element group 544: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1113_sample_completed_
      -- 
    ack_2317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 544_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1113_inst_ack_0, ack => zeropad_CP_182_elements(544)); -- 
    -- CP-element group 545:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 545: predecessors 
    -- CP-element group 545: 	543 
    -- CP-element group 545: successors 
    -- CP-element group 545: 	569 
    -- CP-element group 545: marked-successors 
    -- CP-element group 545: 	305 
    -- CP-element group 545: 	543 
    -- CP-element group 545:  members (3) 
      -- CP-element group 545: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1113_update_completed_
      -- CP-element group 545: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1113_complete/ack
      -- CP-element group 545: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1113_complete/$exit
      -- 
    ack_2322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 545_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1113_inst_ack_1, ack => zeropad_CP_182_elements(545)); -- 
    -- CP-element group 546:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 546: predecessors 
    -- CP-element group 546: 	445 
    -- CP-element group 546: 	453 
    -- CP-element group 546: 	457 
    -- CP-element group 546: 	489 
    -- CP-element group 546: marked-predecessors 
    -- CP-element group 546: 	548 
    -- CP-element group 546: successors 
    -- CP-element group 546: 	548 
    -- CP-element group 546:  members (3) 
      -- CP-element group 546: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1124_Sample/req
      -- CP-element group 546: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1124_Sample/$entry
      -- CP-element group 546: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1124_sample_start_
      -- 
    req_2330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(546), ack => W_condx_xend_ifx_xend238_taken_997_delayed_1_0_1122_inst_req_0); -- 
    zeropad_cp_element_group_546: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_546"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(445) & zeropad_CP_182_elements(453) & zeropad_CP_182_elements(457) & zeropad_CP_182_elements(489) & zeropad_CP_182_elements(548);
      gj_zeropad_cp_element_group_546 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(546), clk => clk, reset => reset); --
    end block;
    -- CP-element group 547:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 547: predecessors 
    -- CP-element group 547: 	115 
    -- CP-element group 547: marked-predecessors 
    -- CP-element group 547: 	549 
    -- CP-element group 547: successors 
    -- CP-element group 547: 	549 
    -- CP-element group 547:  members (3) 
      -- CP-element group 547: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1124_Update/req
      -- CP-element group 547: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1124_Update/$entry
      -- CP-element group 547: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1124_update_start_
      -- 
    req_2335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(547), ack => W_condx_xend_ifx_xend238_taken_997_delayed_1_0_1122_inst_req_1); -- 
    zeropad_cp_element_group_547: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_547"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(549);
      gj_zeropad_cp_element_group_547 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(547), clk => clk, reset => reset); --
    end block;
    -- CP-element group 548:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 548: predecessors 
    -- CP-element group 548: 	546 
    -- CP-element group 548: successors 
    -- CP-element group 548: marked-successors 
    -- CP-element group 548: 	443 
    -- CP-element group 548: 	451 
    -- CP-element group 548: 	455 
    -- CP-element group 548: 	487 
    -- CP-element group 548: 	546 
    -- CP-element group 548:  members (3) 
      -- CP-element group 548: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1124_Sample/ack
      -- CP-element group 548: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1124_Sample/$exit
      -- CP-element group 548: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1124_sample_completed_
      -- 
    ack_2331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 548_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_condx_xend_ifx_xend238_taken_997_delayed_1_0_1122_inst_ack_0, ack => zeropad_CP_182_elements(548)); -- 
    -- CP-element group 549:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 549: predecessors 
    -- CP-element group 549: 	547 
    -- CP-element group 549: successors 
    -- CP-element group 549: 	611 
    -- CP-element group 549: marked-successors 
    -- CP-element group 549: 	137 
    -- CP-element group 549: 	547 
    -- CP-element group 549:  members (3) 
      -- CP-element group 549: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1124_Update/ack
      -- CP-element group 549: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1124_Update/$exit
      -- CP-element group 549: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1124_update_completed_
      -- 
    ack_2336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 549_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_condx_xend_ifx_xend238_taken_997_delayed_1_0_1122_inst_ack_1, ack => zeropad_CP_182_elements(549)); -- 
    -- CP-element group 550:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 550: predecessors 
    -- CP-element group 550: 	142 
    -- CP-element group 550: 	163 
    -- CP-element group 550: marked-predecessors 
    -- CP-element group 550: 	552 
    -- CP-element group 550: successors 
    -- CP-element group 550: 	552 
    -- CP-element group 550:  members (3) 
      -- CP-element group 550: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1131_start/$entry
      -- CP-element group 550: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1131_start/req
      -- CP-element group 550: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1131_sample_start_
      -- 
    req_2344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(550), ack => MUX_1131_inst_req_0); -- 
    zeropad_cp_element_group_550: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_550"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(142) & zeropad_CP_182_elements(163) & zeropad_CP_182_elements(552);
      gj_zeropad_cp_element_group_550 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(550), clk => clk, reset => reset); --
    end block;
    -- CP-element group 551:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 551: predecessors 
    -- CP-element group 551: 	115 
    -- CP-element group 551: marked-predecessors 
    -- CP-element group 551: 	553 
    -- CP-element group 551: successors 
    -- CP-element group 551: 	553 
    -- CP-element group 551:  members (3) 
      -- CP-element group 551: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1131_complete/$entry
      -- CP-element group 551: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1131_complete/req
      -- CP-element group 551: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1131_update_start_
      -- 
    req_2349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(551), ack => MUX_1131_inst_req_1); -- 
    zeropad_cp_element_group_551: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_551"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(553);
      gj_zeropad_cp_element_group_551 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(551), clk => clk, reset => reset); --
    end block;
    -- CP-element group 552:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 552: predecessors 
    -- CP-element group 552: 	550 
    -- CP-element group 552: successors 
    -- CP-element group 552: marked-successors 
    -- CP-element group 552: 	138 
    -- CP-element group 552: 	159 
    -- CP-element group 552: 	550 
    -- CP-element group 552:  members (3) 
      -- CP-element group 552: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1131_start/ack
      -- CP-element group 552: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1131_start/$exit
      -- CP-element group 552: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1131_sample_completed_
      -- 
    ack_2345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 552_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1131_inst_ack_0, ack => zeropad_CP_182_elements(552)); -- 
    -- CP-element group 553:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 553: predecessors 
    -- CP-element group 553: 	551 
    -- CP-element group 553: successors 
    -- CP-element group 553: 	611 
    -- CP-element group 553: marked-successors 
    -- CP-element group 553: 	137 
    -- CP-element group 553: 	551 
    -- CP-element group 553:  members (3) 
      -- CP-element group 553: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1131_update_completed_
      -- CP-element group 553: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1131_complete/$exit
      -- CP-element group 553: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/MUX_1131_complete/ack
      -- 
    ack_2350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 553_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_1131_inst_ack_1, ack => zeropad_CP_182_elements(553)); -- 
    -- CP-element group 554:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 554: predecessors 
    -- CP-element group 554: 	163 
    -- CP-element group 554: marked-predecessors 
    -- CP-element group 554: 	556 
    -- CP-element group 554: successors 
    -- CP-element group 554: 	556 
    -- CP-element group 554:  members (3) 
      -- CP-element group 554: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1142_sample_start_
      -- CP-element group 554: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1142_Sample/$entry
      -- CP-element group 554: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1142_Sample/req
      -- 
    req_2358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(554), ack => W_iNsTr_28_1010_delayed_2_0_1140_inst_req_0); -- 
    zeropad_cp_element_group_554: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_554"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(163) & zeropad_CP_182_elements(556);
      gj_zeropad_cp_element_group_554 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(554), clk => clk, reset => reset); --
    end block;
    -- CP-element group 555:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 555: predecessors 
    -- CP-element group 555: 	115 
    -- CP-element group 555: marked-predecessors 
    -- CP-element group 555: 	557 
    -- CP-element group 555: successors 
    -- CP-element group 555: 	557 
    -- CP-element group 555:  members (3) 
      -- CP-element group 555: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1142_update_start_
      -- CP-element group 555: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1142_Update/$entry
      -- CP-element group 555: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1142_Update/req
      -- 
    req_2363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(555), ack => W_iNsTr_28_1010_delayed_2_0_1140_inst_req_1); -- 
    zeropad_cp_element_group_555: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_555"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(557);
      gj_zeropad_cp_element_group_555 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(555), clk => clk, reset => reset); --
    end block;
    -- CP-element group 556:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 556: predecessors 
    -- CP-element group 556: 	554 
    -- CP-element group 556: successors 
    -- CP-element group 556: marked-successors 
    -- CP-element group 556: 	159 
    -- CP-element group 556: 	554 
    -- CP-element group 556:  members (3) 
      -- CP-element group 556: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1142_sample_completed_
      -- CP-element group 556: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1142_Sample/$exit
      -- CP-element group 556: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1142_Sample/ack
      -- 
    ack_2359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 556_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iNsTr_28_1010_delayed_2_0_1140_inst_ack_0, ack => zeropad_CP_182_elements(556)); -- 
    -- CP-element group 557:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 557: predecessors 
    -- CP-element group 557: 	555 
    -- CP-element group 557: successors 
    -- CP-element group 557: 	611 
    -- CP-element group 557: marked-successors 
    -- CP-element group 557: 	158 
    -- CP-element group 557: 	555 
    -- CP-element group 557:  members (3) 
      -- CP-element group 557: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1142_update_completed_
      -- CP-element group 557: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1142_Update/$exit
      -- CP-element group 557: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1142_Update/ack
      -- 
    ack_2364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 557_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_iNsTr_28_1010_delayed_2_0_1140_inst_ack_1, ack => zeropad_CP_182_elements(557)); -- 
    -- CP-element group 558:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 558: predecessors 
    -- CP-element group 558: 	205 
    -- CP-element group 558: marked-predecessors 
    -- CP-element group 558: 	560 
    -- CP-element group 558: successors 
    -- CP-element group 558: 	560 
    -- CP-element group 558:  members (3) 
      -- CP-element group 558: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1152_Sample/req
      -- CP-element group 558: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1152_Sample/$entry
      -- CP-element group 558: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1152_sample_start_
      -- 
    req_2372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(558), ack => W_output_byte_countx_x0_1017_delayed_2_0_1150_inst_req_0); -- 
    zeropad_cp_element_group_558: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_558"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(205) & zeropad_CP_182_elements(560);
      gj_zeropad_cp_element_group_558 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(558), clk => clk, reset => reset); --
    end block;
    -- CP-element group 559:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 559: predecessors 
    -- CP-element group 559: 	115 
    -- CP-element group 559: marked-predecessors 
    -- CP-element group 559: 	561 
    -- CP-element group 559: successors 
    -- CP-element group 559: 	561 
    -- CP-element group 559:  members (3) 
      -- CP-element group 559: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1152_Update/$entry
      -- CP-element group 559: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1152_update_start_
      -- CP-element group 559: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1152_Update/req
      -- 
    req_2377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(559), ack => W_output_byte_countx_x0_1017_delayed_2_0_1150_inst_req_1); -- 
    zeropad_cp_element_group_559: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_559"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(561);
      gj_zeropad_cp_element_group_559 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(559), clk => clk, reset => reset); --
    end block;
    -- CP-element group 560:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 560: predecessors 
    -- CP-element group 560: 	558 
    -- CP-element group 560: successors 
    -- CP-element group 560: marked-successors 
    -- CP-element group 560: 	201 
    -- CP-element group 560: 	558 
    -- CP-element group 560:  members (3) 
      -- CP-element group 560: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1152_Sample/ack
      -- CP-element group 560: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1152_Sample/$exit
      -- CP-element group 560: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1152_sample_completed_
      -- 
    ack_2373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 560_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_byte_countx_x0_1017_delayed_2_0_1150_inst_ack_0, ack => zeropad_CP_182_elements(560)); -- 
    -- CP-element group 561:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 561: predecessors 
    -- CP-element group 561: 	559 
    -- CP-element group 561: successors 
    -- CP-element group 561: 	611 
    -- CP-element group 561: marked-successors 
    -- CP-element group 561: 	179 
    -- CP-element group 561: 	200 
    -- CP-element group 561: 	305 
    -- CP-element group 561: 	559 
    -- CP-element group 561:  members (3) 
      -- CP-element group 561: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1152_Update/$exit
      -- CP-element group 561: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1152_update_completed_
      -- CP-element group 561: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1152_Update/ack
      -- 
    ack_2378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 561_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_byte_countx_x0_1017_delayed_2_0_1150_inst_ack_1, ack => zeropad_CP_182_elements(561)); -- 
    -- CP-element group 562:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 562: predecessors 
    -- CP-element group 562: 	566 
    -- CP-element group 562: marked-predecessors 
    -- CP-element group 562: 	567 
    -- CP-element group 562: successors 
    -- CP-element group 562: 	567 
    -- CP-element group 562:  members (3) 
      -- CP-element group 562: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_1188_request/$entry
      -- CP-element group 562: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_1188_request/req
      -- CP-element group 562: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_1188_sample_start_
      -- 
    req_2418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(562), ack => addr_of_1188_final_reg_req_0); -- 
    zeropad_cp_element_group_562: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_562"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(566) & zeropad_CP_182_elements(567);
      gj_zeropad_cp_element_group_562 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(562), clk => clk, reset => reset); --
    end block;
    -- CP-element group 563:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 563: predecessors 
    -- CP-element group 563: 	112 
    -- CP-element group 563: marked-predecessors 
    -- CP-element group 563: 	568 
    -- CP-element group 563: 	571 
    -- CP-element group 563: successors 
    -- CP-element group 563: 	568 
    -- CP-element group 563:  members (3) 
      -- CP-element group 563: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_1188_complete/$entry
      -- CP-element group 563: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_1188_complete/req
      -- CP-element group 563: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_1188_update_start_
      -- 
    req_2423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(563), ack => addr_of_1188_final_reg_req_1); -- 
    zeropad_cp_element_group_563: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_563"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(568) & zeropad_CP_182_elements(571);
      gj_zeropad_cp_element_group_563 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(563), clk => clk, reset => reset); --
    end block;
    -- CP-element group 564:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 564: predecessors 
    -- CP-element group 564: 	112 
    -- CP-element group 564: marked-predecessors 
    -- CP-element group 564: 	566 
    -- CP-element group 564: 	567 
    -- CP-element group 564: successors 
    -- CP-element group 564: 	566 
    -- CP-element group 564:  members (3) 
      -- CP-element group 564: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_final_index_sum_regn_Update/req
      -- CP-element group 564: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_final_index_sum_regn_Update/$entry
      -- CP-element group 564: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_final_index_sum_regn_update_start
      -- 
    req_2408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(564), ack => array_obj_ref_1187_index_offset_req_1); -- 
    zeropad_cp_element_group_564: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_564"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(566) & zeropad_CP_182_elements(567);
      gj_zeropad_cp_element_group_564 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(564), clk => clk, reset => reset); --
    end block;
    -- CP-element group 565:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 565: predecessors 
    -- CP-element group 565: 	184 
    -- CP-element group 565: successors 
    -- CP-element group 565: 	611 
    -- CP-element group 565: marked-successors 
    -- CP-element group 565: 	180 
    -- CP-element group 565:  members (3) 
      -- CP-element group 565: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_final_index_sum_regn_Sample/ack
      -- CP-element group 565: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_final_index_sum_regn_Sample/$exit
      -- CP-element group 565: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_final_index_sum_regn_sample_complete
      -- 
    ack_2404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 565_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1187_index_offset_ack_0, ack => zeropad_CP_182_elements(565)); -- 
    -- CP-element group 566:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 566: predecessors 
    -- CP-element group 566: 	564 
    -- CP-element group 566: successors 
    -- CP-element group 566: 	562 
    -- CP-element group 566: marked-successors 
    -- CP-element group 566: 	564 
    -- CP-element group 566:  members (8) 
      -- CP-element group 566: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_final_index_sum_regn_Update/ack
      -- CP-element group 566: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_base_plus_offset/$entry
      -- CP-element group 566: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_base_plus_offset/sum_rename_req
      -- CP-element group 566: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_base_plus_offset/$exit
      -- CP-element group 566: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_base_plus_offset/sum_rename_ack
      -- CP-element group 566: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_final_index_sum_regn_Update/$exit
      -- CP-element group 566: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_offset_calculated
      -- CP-element group 566: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/array_obj_ref_1187_root_address_calculated
      -- 
    ack_2409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 566_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1187_index_offset_ack_1, ack => zeropad_CP_182_elements(566)); -- 
    -- CP-element group 567:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 567: predecessors 
    -- CP-element group 567: 	562 
    -- CP-element group 567: successors 
    -- CP-element group 567: marked-successors 
    -- CP-element group 567: 	562 
    -- CP-element group 567: 	564 
    -- CP-element group 567:  members (3) 
      -- CP-element group 567: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_1188_request/$exit
      -- CP-element group 567: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_1188_request/ack
      -- CP-element group 567: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_1188_sample_completed_
      -- 
    ack_2419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 567_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1188_final_reg_ack_0, ack => zeropad_CP_182_elements(567)); -- 
    -- CP-element group 568:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 568: predecessors 
    -- CP-element group 568: 	563 
    -- CP-element group 568: successors 
    -- CP-element group 568: 	569 
    -- CP-element group 568: marked-successors 
    -- CP-element group 568: 	563 
    -- CP-element group 568:  members (19) 
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_1188_complete/$exit
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_1188_complete/ack
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_base_address_calculated
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_word_address_calculated
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_root_address_calculated
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_base_address_resized
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_base_addr_resize/$entry
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_base_addr_resize/$exit
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_base_addr_resize/base_resize_req
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_base_addr_resize/base_resize_ack
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_base_plus_offset/$entry
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_base_plus_offset/$exit
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_base_plus_offset/sum_rename_req
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_base_plus_offset/sum_rename_ack
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_word_addrgen/$entry
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_word_addrgen/$exit
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_word_addrgen/root_register_req
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_word_addrgen/root_register_ack
      -- CP-element group 568: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/addr_of_1188_update_completed_
      -- 
    ack_2424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 568_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1188_final_reg_ack_1, ack => zeropad_CP_182_elements(568)); -- 
    -- CP-element group 569:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 569: predecessors 
    -- CP-element group 569: 	366 
    -- CP-element group 569: 	374 
    -- CP-element group 569: 	386 
    -- CP-element group 569: 	445 
    -- CP-element group 569: 	453 
    -- CP-element group 569: 	457 
    -- CP-element group 569: 	489 
    -- CP-element group 569: 	545 
    -- CP-element group 569: 	568 
    -- CP-element group 569: 	610 
    -- CP-element group 569: marked-predecessors 
    -- CP-element group 569: 	571 
    -- CP-element group 569: successors 
    -- CP-element group 569: 	571 
    -- CP-element group 569:  members (9) 
      -- CP-element group 569: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Sample/ptr_deref_1192_Split/$exit
      -- CP-element group 569: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Sample/word_access_start/word_0/$entry
      -- CP-element group 569: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Sample/word_access_start/word_0/rr
      -- CP-element group 569: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Sample/ptr_deref_1192_Split/$entry
      -- CP-element group 569: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Sample/ptr_deref_1192_Split/split_ack
      -- CP-element group 569: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Sample/word_access_start/$entry
      -- CP-element group 569: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Sample/ptr_deref_1192_Split/split_req
      -- CP-element group 569: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_sample_start_
      -- CP-element group 569: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Sample/$entry
      -- 
    rr_2462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(569), ack => ptr_deref_1192_store_0_req_0); -- 
    zeropad_cp_element_group_569: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 1);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_569"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(366) & zeropad_CP_182_elements(374) & zeropad_CP_182_elements(386) & zeropad_CP_182_elements(445) & zeropad_CP_182_elements(453) & zeropad_CP_182_elements(457) & zeropad_CP_182_elements(489) & zeropad_CP_182_elements(545) & zeropad_CP_182_elements(568) & zeropad_CP_182_elements(610) & zeropad_CP_182_elements(571);
      gj_zeropad_cp_element_group_569 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(569), clk => clk, reset => reset); --
    end block;
    -- CP-element group 570:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 570: predecessors 
    -- CP-element group 570: marked-predecessors 
    -- CP-element group 570: 	572 
    -- CP-element group 570: successors 
    -- CP-element group 570: 	572 
    -- CP-element group 570:  members (5) 
      -- CP-element group 570: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Update/word_access_complete/word_0/$entry
      -- CP-element group 570: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Update/$entry
      -- CP-element group 570: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Update/word_access_complete/$entry
      -- CP-element group 570: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_update_start_
      -- CP-element group 570: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Update/word_access_complete/word_0/cr
      -- 
    cr_2473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(570), ack => ptr_deref_1192_store_0_req_1); -- 
    zeropad_cp_element_group_570: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_570"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad_CP_182_elements(572);
      gj_zeropad_cp_element_group_570 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(570), clk => clk, reset => reset); --
    end block;
    -- CP-element group 571:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 571: predecessors 
    -- CP-element group 571: 	569 
    -- CP-element group 571: successors 
    -- CP-element group 571: 	611 
    -- CP-element group 571: marked-successors 
    -- CP-element group 571: 	364 
    -- CP-element group 571: 	372 
    -- CP-element group 571: 	384 
    -- CP-element group 571: 	398 
    -- CP-element group 571: 	443 
    -- CP-element group 571: 	451 
    -- CP-element group 571: 	455 
    -- CP-element group 571: 	487 
    -- CP-element group 571: 	543 
    -- CP-element group 571: 	563 
    -- CP-element group 571: 	569 
    -- CP-element group 571:  members (6) 
      -- CP-element group 571: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Sample/word_access_start/word_0/ra
      -- CP-element group 571: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Sample/word_access_start/$exit
      -- CP-element group 571: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Sample/word_access_start/word_0/$exit
      -- CP-element group 571: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Sample/$exit
      -- CP-element group 571: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_sample_completed_
      -- CP-element group 571: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ring_reenable_memory_space_0
      -- 
    ra_2463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 571_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1192_store_0_ack_0, ack => zeropad_CP_182_elements(571)); -- 
    -- CP-element group 572:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 572: predecessors 
    -- CP-element group 572: 	570 
    -- CP-element group 572: successors 
    -- CP-element group 572: 	611 
    -- CP-element group 572: marked-successors 
    -- CP-element group 572: 	570 
    -- CP-element group 572:  members (5) 
      -- CP-element group 572: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Update/$exit
      -- CP-element group 572: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Update/word_access_complete/$exit
      -- CP-element group 572: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_update_completed_
      -- CP-element group 572: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Update/word_access_complete/word_0/$exit
      -- CP-element group 572: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_1192_Update/word_access_complete/word_0/ca
      -- 
    ca_2474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 572_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1192_store_0_ack_1, ack => zeropad_CP_182_elements(572)); -- 
    -- CP-element group 573:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 573: predecessors 
    -- CP-element group 573: 	184 
    -- CP-element group 573: marked-predecessors 
    -- CP-element group 573: 	575 
    -- CP-element group 573: successors 
    -- CP-element group 573: 	575 
    -- CP-element group 573:  members (3) 
      -- CP-element group 573: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1197_Sample/req
      -- CP-element group 573: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1197_Sample/$entry
      -- CP-element group 573: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1197_sample_start_
      -- 
    req_2482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(573), ack => W_add_outx_x1_1059_delayed_2_0_1195_inst_req_0); -- 
    zeropad_cp_element_group_573: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_573"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(184) & zeropad_CP_182_elements(575);
      gj_zeropad_cp_element_group_573 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(573), clk => clk, reset => reset); --
    end block;
    -- CP-element group 574:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 574: predecessors 
    -- CP-element group 574: 	115 
    -- CP-element group 574: marked-predecessors 
    -- CP-element group 574: 	576 
    -- CP-element group 574: successors 
    -- CP-element group 574: 	576 
    -- CP-element group 574:  members (3) 
      -- CP-element group 574: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1197_Update/req
      -- CP-element group 574: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1197_Update/$entry
      -- CP-element group 574: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1197_update_start_
      -- 
    req_2487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(574), ack => W_add_outx_x1_1059_delayed_2_0_1195_inst_req_1); -- 
    zeropad_cp_element_group_574: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_574"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(576);
      gj_zeropad_cp_element_group_574 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(574), clk => clk, reset => reset); --
    end block;
    -- CP-element group 575:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 575: predecessors 
    -- CP-element group 575: 	573 
    -- CP-element group 575: successors 
    -- CP-element group 575: marked-successors 
    -- CP-element group 575: 	180 
    -- CP-element group 575: 	573 
    -- CP-element group 575:  members (3) 
      -- CP-element group 575: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1197_Sample/ack
      -- CP-element group 575: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1197_Sample/$exit
      -- CP-element group 575: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1197_sample_completed_
      -- 
    ack_2483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 575_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_outx_x1_1059_delayed_2_0_1195_inst_ack_0, ack => zeropad_CP_182_elements(575)); -- 
    -- CP-element group 576:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 576: predecessors 
    -- CP-element group 576: 	574 
    -- CP-element group 576: successors 
    -- CP-element group 576: 	611 
    -- CP-element group 576: marked-successors 
    -- CP-element group 576: 	179 
    -- CP-element group 576: 	574 
    -- CP-element group 576:  members (3) 
      -- CP-element group 576: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1197_Update/ack
      -- CP-element group 576: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1197_Update/$exit
      -- CP-element group 576: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1197_update_completed_
      -- 
    ack_2488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 576_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_outx_x1_1059_delayed_2_0_1195_inst_ack_1, ack => zeropad_CP_182_elements(576)); -- 
    -- CP-element group 577:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 577: predecessors 
    -- CP-element group 577: 	184 
    -- CP-element group 577: marked-predecessors 
    -- CP-element group 577: 	579 
    -- CP-element group 577: successors 
    -- CP-element group 577: 	579 
    -- CP-element group 577:  members (3) 
      -- CP-element group 577: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1210_Sample/rr
      -- CP-element group 577: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1210_Sample/$entry
      -- CP-element group 577: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1210_sample_start_
      -- 
    rr_2496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(577), ack => type_cast_1210_inst_req_0); -- 
    zeropad_cp_element_group_577: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_577"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(184) & zeropad_CP_182_elements(579);
      gj_zeropad_cp_element_group_577 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(577), clk => clk, reset => reset); --
    end block;
    -- CP-element group 578:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 578: predecessors 
    -- CP-element group 578: 	115 
    -- CP-element group 578: marked-predecessors 
    -- CP-element group 578: 	580 
    -- CP-element group 578: successors 
    -- CP-element group 578: 	580 
    -- CP-element group 578:  members (3) 
      -- CP-element group 578: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1210_Update/$entry
      -- CP-element group 578: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1210_Update/cr
      -- CP-element group 578: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1210_update_start_
      -- 
    cr_2501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(578), ack => type_cast_1210_inst_req_1); -- 
    zeropad_cp_element_group_578: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_578"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(580);
      gj_zeropad_cp_element_group_578 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(578), clk => clk, reset => reset); --
    end block;
    -- CP-element group 579:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 579: predecessors 
    -- CP-element group 579: 	577 
    -- CP-element group 579: successors 
    -- CP-element group 579: marked-successors 
    -- CP-element group 579: 	180 
    -- CP-element group 579: 	577 
    -- CP-element group 579:  members (3) 
      -- CP-element group 579: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1210_Sample/ra
      -- CP-element group 579: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1210_Sample/$exit
      -- CP-element group 579: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1210_sample_completed_
      -- 
    ra_2497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 579_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1210_inst_ack_0, ack => zeropad_CP_182_elements(579)); -- 
    -- CP-element group 580:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 580: predecessors 
    -- CP-element group 580: 	578 
    -- CP-element group 580: successors 
    -- CP-element group 580: 	611 
    -- CP-element group 580: marked-successors 
    -- CP-element group 580: 	179 
    -- CP-element group 580: 	578 
    -- CP-element group 580:  members (3) 
      -- CP-element group 580: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1210_Update/ca
      -- CP-element group 580: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1210_Update/$exit
      -- CP-element group 580: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1210_update_completed_
      -- 
    ca_2502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 580_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1210_inst_ack_1, ack => zeropad_CP_182_elements(580)); -- 
    -- CP-element group 581:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 581: predecessors 
    -- CP-element group 581: 	289 
    -- CP-element group 581: marked-predecessors 
    -- CP-element group 581: 	583 
    -- CP-element group 581: successors 
    -- CP-element group 581: 	583 
    -- CP-element group 581:  members (3) 
      -- CP-element group 581: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1251_sample_start_
      -- CP-element group 581: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1251_Sample/$entry
      -- CP-element group 581: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1251_Sample/rr
      -- 
    rr_2510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(581), ack => type_cast_1251_inst_req_0); -- 
    zeropad_cp_element_group_581: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_581"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(289) & zeropad_CP_182_elements(583);
      gj_zeropad_cp_element_group_581 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(581), clk => clk, reset => reset); --
    end block;
    -- CP-element group 582:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 582: predecessors 
    -- CP-element group 582: 	115 
    -- CP-element group 582: marked-predecessors 
    -- CP-element group 582: 	584 
    -- CP-element group 582: 	591 
    -- CP-element group 582: successors 
    -- CP-element group 582: 	584 
    -- CP-element group 582:  members (3) 
      -- CP-element group 582: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1251_update_start_
      -- CP-element group 582: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1251_Update/$entry
      -- CP-element group 582: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1251_Update/cr
      -- 
    cr_2515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(582), ack => type_cast_1251_inst_req_1); -- 
    zeropad_cp_element_group_582: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_582"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(584) & zeropad_CP_182_elements(591);
      gj_zeropad_cp_element_group_582 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(582), clk => clk, reset => reset); --
    end block;
    -- CP-element group 583:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 583: predecessors 
    -- CP-element group 583: 	581 
    -- CP-element group 583: successors 
    -- CP-element group 583: marked-successors 
    -- CP-element group 583: 	285 
    -- CP-element group 583: 	581 
    -- CP-element group 583:  members (3) 
      -- CP-element group 583: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1251_sample_completed_
      -- CP-element group 583: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1251_Sample/$exit
      -- CP-element group 583: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1251_Sample/ra
      -- 
    ra_2511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 583_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1251_inst_ack_0, ack => zeropad_CP_182_elements(583)); -- 
    -- CP-element group 584:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 584: predecessors 
    -- CP-element group 584: 	582 
    -- CP-element group 584: successors 
    -- CP-element group 584: 	589 
    -- CP-element group 584: marked-successors 
    -- CP-element group 584: 	284 
    -- CP-element group 584: 	582 
    -- CP-element group 584:  members (3) 
      -- CP-element group 584: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1251_update_completed_
      -- CP-element group 584: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1251_Update/$exit
      -- CP-element group 584: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1251_Update/ca
      -- 
    ca_2516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 584_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1251_inst_ack_1, ack => zeropad_CP_182_elements(584)); -- 
    -- CP-element group 585:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 585: predecessors 
    -- CP-element group 585: 	112 
    -- CP-element group 585: marked-predecessors 
    -- CP-element group 585: 	587 
    -- CP-element group 585: successors 
    -- CP-element group 585: 	587 
    -- CP-element group 585:  members (3) 
      -- CP-element group 585: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1255_sample_start_
      -- CP-element group 585: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1255_Sample/$entry
      -- CP-element group 585: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1255_Sample/rr
      -- 
    rr_2524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(585), ack => type_cast_1255_inst_req_0); -- 
    zeropad_cp_element_group_585: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_585"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(112) & zeropad_CP_182_elements(587);
      gj_zeropad_cp_element_group_585 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(585), clk => clk, reset => reset); --
    end block;
    -- CP-element group 586:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 586: predecessors 
    -- CP-element group 586: 	115 
    -- CP-element group 586: marked-predecessors 
    -- CP-element group 586: 	588 
    -- CP-element group 586: 	591 
    -- CP-element group 586: successors 
    -- CP-element group 586: 	588 
    -- CP-element group 586:  members (3) 
      -- CP-element group 586: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1255_update_start_
      -- CP-element group 586: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1255_Update/$entry
      -- CP-element group 586: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1255_Update/cr
      -- 
    cr_2529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(586), ack => type_cast_1255_inst_req_1); -- 
    zeropad_cp_element_group_586: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_586"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(588) & zeropad_CP_182_elements(591);
      gj_zeropad_cp_element_group_586 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(586), clk => clk, reset => reset); --
    end block;
    -- CP-element group 587:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 587: predecessors 
    -- CP-element group 587: 	585 
    -- CP-element group 587: successors 
    -- CP-element group 587: marked-successors 
    -- CP-element group 587: 	585 
    -- CP-element group 587:  members (3) 
      -- CP-element group 587: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1255_sample_completed_
      -- CP-element group 587: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1255_Sample/$exit
      -- CP-element group 587: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1255_Sample/ra
      -- 
    ra_2525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 587_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1255_inst_ack_0, ack => zeropad_CP_182_elements(587)); -- 
    -- CP-element group 588:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 588: predecessors 
    -- CP-element group 588: 	586 
    -- CP-element group 588: successors 
    -- CP-element group 588: 	589 
    -- CP-element group 588: marked-successors 
    -- CP-element group 588: 	284 
    -- CP-element group 588: 	586 
    -- CP-element group 588:  members (3) 
      -- CP-element group 588: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1255_update_completed_
      -- CP-element group 588: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1255_Update/$exit
      -- CP-element group 588: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1255_Update/ca
      -- 
    ca_2530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 588_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1255_inst_ack_1, ack => zeropad_CP_182_elements(588)); -- 
    -- CP-element group 589:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 589: predecessors 
    -- CP-element group 589: 	584 
    -- CP-element group 589: 	588 
    -- CP-element group 589: marked-predecessors 
    -- CP-element group 589: 	591 
    -- CP-element group 589: successors 
    -- CP-element group 589: 	591 
    -- CP-element group 589:  members (3) 
      -- CP-element group 589: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1271_sample_start_
      -- CP-element group 589: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1271_Sample/$entry
      -- CP-element group 589: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1271_Sample/rr
      -- 
    rr_2538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(589), ack => type_cast_1271_inst_req_0); -- 
    zeropad_cp_element_group_589: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_589"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(584) & zeropad_CP_182_elements(588) & zeropad_CP_182_elements(591);
      gj_zeropad_cp_element_group_589 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(589), clk => clk, reset => reset); --
    end block;
    -- CP-element group 590:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 590: predecessors 
    -- CP-element group 590: 	115 
    -- CP-element group 590: marked-predecessors 
    -- CP-element group 590: 	592 
    -- CP-element group 590: 	603 
    -- CP-element group 590: successors 
    -- CP-element group 590: 	592 
    -- CP-element group 590:  members (3) 
      -- CP-element group 590: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1271_update_start_
      -- CP-element group 590: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1271_Update/$entry
      -- CP-element group 590: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1271_Update/cr
      -- 
    cr_2543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(590), ack => type_cast_1271_inst_req_1); -- 
    zeropad_cp_element_group_590: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_590"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(592) & zeropad_CP_182_elements(603);
      gj_zeropad_cp_element_group_590 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(590), clk => clk, reset => reset); --
    end block;
    -- CP-element group 591:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 591: predecessors 
    -- CP-element group 591: 	589 
    -- CP-element group 591: successors 
    -- CP-element group 591: marked-successors 
    -- CP-element group 591: 	582 
    -- CP-element group 591: 	586 
    -- CP-element group 591: 	589 
    -- CP-element group 591:  members (3) 
      -- CP-element group 591: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1271_sample_completed_
      -- CP-element group 591: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1271_Sample/$exit
      -- CP-element group 591: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1271_Sample/ra
      -- 
    ra_2539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 591_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1271_inst_ack_0, ack => zeropad_CP_182_elements(591)); -- 
    -- CP-element group 592:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 592: predecessors 
    -- CP-element group 592: 	590 
    -- CP-element group 592: successors 
    -- CP-element group 592: 	601 
    -- CP-element group 592: marked-successors 
    -- CP-element group 592: 	263 
    -- CP-element group 592: 	590 
    -- CP-element group 592:  members (3) 
      -- CP-element group 592: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1271_update_completed_
      -- CP-element group 592: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1271_Update/$exit
      -- CP-element group 592: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1271_Update/ca
      -- 
    ca_2544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 592_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1271_inst_ack_1, ack => zeropad_CP_182_elements(592)); -- 
    -- CP-element group 593:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 593: predecessors 
    -- CP-element group 593: 	268 
    -- CP-element group 593: marked-predecessors 
    -- CP-element group 593: 	595 
    -- CP-element group 593: successors 
    -- CP-element group 593: 	595 
    -- CP-element group 593:  members (3) 
      -- CP-element group 593: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1281_sample_start_
      -- CP-element group 593: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1281_Sample/$entry
      -- CP-element group 593: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1281_Sample/req
      -- 
    req_2552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(593), ack => W_o1x_x1_1134_delayed_2_0_1279_inst_req_0); -- 
    zeropad_cp_element_group_593: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_593"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(268) & zeropad_CP_182_elements(595);
      gj_zeropad_cp_element_group_593 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(593), clk => clk, reset => reset); --
    end block;
    -- CP-element group 594:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 594: predecessors 
    -- CP-element group 594: 	115 
    -- CP-element group 594: marked-predecessors 
    -- CP-element group 594: 	596 
    -- CP-element group 594: 	603 
    -- CP-element group 594: successors 
    -- CP-element group 594: 	596 
    -- CP-element group 594:  members (3) 
      -- CP-element group 594: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1281_update_start_
      -- CP-element group 594: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1281_Update/$entry
      -- CP-element group 594: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1281_Update/req
      -- 
    req_2557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(594), ack => W_o1x_x1_1134_delayed_2_0_1279_inst_req_1); -- 
    zeropad_cp_element_group_594: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_594"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(596) & zeropad_CP_182_elements(603);
      gj_zeropad_cp_element_group_594 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(594), clk => clk, reset => reset); --
    end block;
    -- CP-element group 595:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 595: predecessors 
    -- CP-element group 595: 	593 
    -- CP-element group 595: successors 
    -- CP-element group 595: marked-successors 
    -- CP-element group 595: 	264 
    -- CP-element group 595: 	593 
    -- CP-element group 595:  members (3) 
      -- CP-element group 595: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1281_sample_completed_
      -- CP-element group 595: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1281_Sample/$exit
      -- CP-element group 595: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1281_Sample/ack
      -- 
    ack_2553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 595_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_o1x_x1_1134_delayed_2_0_1279_inst_ack_0, ack => zeropad_CP_182_elements(595)); -- 
    -- CP-element group 596:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 596: predecessors 
    -- CP-element group 596: 	594 
    -- CP-element group 596: successors 
    -- CP-element group 596: 	601 
    -- CP-element group 596: marked-successors 
    -- CP-element group 596: 	263 
    -- CP-element group 596: 	594 
    -- CP-element group 596:  members (3) 
      -- CP-element group 596: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1281_update_completed_
      -- CP-element group 596: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1281_Update/$exit
      -- CP-element group 596: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1281_Update/ack
      -- 
    ack_2558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 596_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_o1x_x1_1134_delayed_2_0_1279_inst_ack_1, ack => zeropad_CP_182_elements(596)); -- 
    -- CP-element group 597:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 597: predecessors 
    -- CP-element group 597: 	289 
    -- CP-element group 597: marked-predecessors 
    -- CP-element group 597: 	599 
    -- CP-element group 597: successors 
    -- CP-element group 597: 	599 
    -- CP-element group 597:  members (3) 
      -- CP-element group 597: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1289_sample_start_
      -- CP-element group 597: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1289_Sample/$entry
      -- CP-element group 597: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1289_Sample/req
      -- 
    req_2566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(597), ack => W_inc265_1139_delayed_1_0_1287_inst_req_0); -- 
    zeropad_cp_element_group_597: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_597"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(289) & zeropad_CP_182_elements(599);
      gj_zeropad_cp_element_group_597 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(597), clk => clk, reset => reset); --
    end block;
    -- CP-element group 598:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 598: predecessors 
    -- CP-element group 598: 	115 
    -- CP-element group 598: marked-predecessors 
    -- CP-element group 598: 	600 
    -- CP-element group 598: successors 
    -- CP-element group 598: 	600 
    -- CP-element group 598:  members (3) 
      -- CP-element group 598: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1289_update_start_
      -- CP-element group 598: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1289_Update/$entry
      -- CP-element group 598: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1289_Update/req
      -- 
    req_2571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(598), ack => W_inc265_1139_delayed_1_0_1287_inst_req_1); -- 
    zeropad_cp_element_group_598: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_598"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(600);
      gj_zeropad_cp_element_group_598 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(598), clk => clk, reset => reset); --
    end block;
    -- CP-element group 599:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 599: predecessors 
    -- CP-element group 599: 	597 
    -- CP-element group 599: successors 
    -- CP-element group 599: marked-successors 
    -- CP-element group 599: 	285 
    -- CP-element group 599: 	597 
    -- CP-element group 599:  members (3) 
      -- CP-element group 599: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1289_sample_completed_
      -- CP-element group 599: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1289_Sample/$exit
      -- CP-element group 599: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1289_Sample/ack
      -- 
    ack_2567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 599_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_inc265_1139_delayed_1_0_1287_inst_ack_0, ack => zeropad_CP_182_elements(599)); -- 
    -- CP-element group 600:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 600: predecessors 
    -- CP-element group 600: 	598 
    -- CP-element group 600: successors 
    -- CP-element group 600: 	611 
    -- CP-element group 600: marked-successors 
    -- CP-element group 600: 	284 
    -- CP-element group 600: 	598 
    -- CP-element group 600:  members (3) 
      -- CP-element group 600: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1289_update_completed_
      -- CP-element group 600: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1289_Update/$exit
      -- CP-element group 600: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1289_Update/ack
      -- 
    ack_2572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 600_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_inc265_1139_delayed_1_0_1287_inst_ack_1, ack => zeropad_CP_182_elements(600)); -- 
    -- CP-element group 601:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 601: predecessors 
    -- CP-element group 601: 	592 
    -- CP-element group 601: 	596 
    -- CP-element group 601: marked-predecessors 
    -- CP-element group 601: 	603 
    -- CP-element group 601: successors 
    -- CP-element group 601: 	603 
    -- CP-element group 601:  members (3) 
      -- CP-element group 601: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1304_sample_start_
      -- CP-element group 601: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1304_Sample/$entry
      -- CP-element group 601: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1304_Sample/rr
      -- 
    rr_2580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(601), ack => type_cast_1304_inst_req_0); -- 
    zeropad_cp_element_group_601: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_601"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(592) & zeropad_CP_182_elements(596) & zeropad_CP_182_elements(603);
      gj_zeropad_cp_element_group_601 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(601), clk => clk, reset => reset); --
    end block;
    -- CP-element group 602:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 602: predecessors 
    -- CP-element group 602: 	115 
    -- CP-element group 602: marked-predecessors 
    -- CP-element group 602: 	604 
    -- CP-element group 602: successors 
    -- CP-element group 602: 	604 
    -- CP-element group 602:  members (3) 
      -- CP-element group 602: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1304_update_start_
      -- CP-element group 602: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1304_Update/$entry
      -- CP-element group 602: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1304_Update/cr
      -- 
    cr_2585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(602), ack => type_cast_1304_inst_req_1); -- 
    zeropad_cp_element_group_602: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_602"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(604);
      gj_zeropad_cp_element_group_602 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(602), clk => clk, reset => reset); --
    end block;
    -- CP-element group 603:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 603: predecessors 
    -- CP-element group 603: 	601 
    -- CP-element group 603: successors 
    -- CP-element group 603: marked-successors 
    -- CP-element group 603: 	590 
    -- CP-element group 603: 	594 
    -- CP-element group 603: 	601 
    -- CP-element group 603:  members (3) 
      -- CP-element group 603: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1304_sample_completed_
      -- CP-element group 603: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1304_Sample/$exit
      -- CP-element group 603: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1304_Sample/ra
      -- 
    ra_2581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 603_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1304_inst_ack_0, ack => zeropad_CP_182_elements(603)); -- 
    -- CP-element group 604:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 604: predecessors 
    -- CP-element group 604: 	602 
    -- CP-element group 604: successors 
    -- CP-element group 604: 	113 
    -- CP-element group 604: marked-successors 
    -- CP-element group 604: 	242 
    -- CP-element group 604: 	602 
    -- CP-element group 604:  members (3) 
      -- CP-element group 604: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1304_update_completed_
      -- CP-element group 604: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1304_Update/$exit
      -- CP-element group 604: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/type_cast_1304_Update/ca
      -- 
    ca_2586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 604_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1304_inst_ack_1, ack => zeropad_CP_182_elements(604)); -- 
    -- CP-element group 605:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 605: predecessors 
    -- CP-element group 605: 	247 
    -- CP-element group 605: marked-predecessors 
    -- CP-element group 605: 	607 
    -- CP-element group 605: successors 
    -- CP-element group 605: 	607 
    -- CP-element group 605:  members (3) 
      -- CP-element group 605: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1308_sample_start_
      -- CP-element group 605: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1308_Sample/$entry
      -- CP-element group 605: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1308_Sample/req
      -- 
    req_2594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(605), ack => W_o0x_x1_1155_delayed_3_0_1306_inst_req_0); -- 
    zeropad_cp_element_group_605: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_605"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(247) & zeropad_CP_182_elements(607);
      gj_zeropad_cp_element_group_605 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(605), clk => clk, reset => reset); --
    end block;
    -- CP-element group 606:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 606: predecessors 
    -- CP-element group 606: 	115 
    -- CP-element group 606: marked-predecessors 
    -- CP-element group 606: 	608 
    -- CP-element group 606: successors 
    -- CP-element group 606: 	608 
    -- CP-element group 606:  members (3) 
      -- CP-element group 606: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1308_update_start_
      -- CP-element group 606: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1308_Update/$entry
      -- CP-element group 606: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1308_Update/req
      -- 
    req_2599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(606), ack => W_o0x_x1_1155_delayed_3_0_1306_inst_req_1); -- 
    zeropad_cp_element_group_606: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_606"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(115) & zeropad_CP_182_elements(608);
      gj_zeropad_cp_element_group_606 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(606), clk => clk, reset => reset); --
    end block;
    -- CP-element group 607:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 607: predecessors 
    -- CP-element group 607: 	605 
    -- CP-element group 607: successors 
    -- CP-element group 607: marked-successors 
    -- CP-element group 607: 	243 
    -- CP-element group 607: 	605 
    -- CP-element group 607:  members (3) 
      -- CP-element group 607: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1308_sample_completed_
      -- CP-element group 607: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1308_Sample/$exit
      -- CP-element group 607: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1308_Sample/ack
      -- 
    ack_2595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 607_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_o0x_x1_1155_delayed_3_0_1306_inst_ack_0, ack => zeropad_CP_182_elements(607)); -- 
    -- CP-element group 608:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 608: predecessors 
    -- CP-element group 608: 	606 
    -- CP-element group 608: successors 
    -- CP-element group 608: 	113 
    -- CP-element group 608: marked-successors 
    -- CP-element group 608: 	242 
    -- CP-element group 608: 	606 
    -- CP-element group 608:  members (3) 
      -- CP-element group 608: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1308_update_completed_
      -- CP-element group 608: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1308_Update/$exit
      -- CP-element group 608: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/assign_stmt_1308_Update/ack
      -- 
    ack_2600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 608_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_o0x_x1_1155_delayed_3_0_1306_inst_ack_1, ack => zeropad_CP_182_elements(608)); -- 
    -- CP-element group 609:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 609: predecessors 
    -- CP-element group 609: 	112 
    -- CP-element group 609: successors 
    -- CP-element group 609: 	113 
    -- CP-element group 609:  members (1) 
      -- CP-element group 609: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group zeropad_CP_182_elements(609) is a control-delay.
    cp_element_609_delay: control_delay_element  generic map(name => " 609_delay", delay_value => 1)  port map(req => zeropad_CP_182_elements(112), ack => zeropad_CP_182_elements(609), clk => clk, reset =>reset);
    -- CP-element group 610:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 610: predecessors 
    -- CP-element group 610: 	400 
    -- CP-element group 610: successors 
    -- CP-element group 610: 	569 
    -- CP-element group 610:  members (1) 
      -- CP-element group 610: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/ptr_deref_798_ptr_deref_1192_delay
      -- 
    -- Element group zeropad_CP_182_elements(610) is a control-delay.
    cp_element_610_delay: control_delay_element  generic map(name => " 610_delay", delay_value => 1)  port map(req => zeropad_CP_182_elements(400), ack => zeropad_CP_182_elements(610), clk => clk, reset =>reset);
    -- CP-element group 611:  join  transition  bypass  pipeline-parent 
    -- CP-element group 611: predecessors 
    -- CP-element group 611: 	354 
    -- CP-element group 611: 	358 
    -- CP-element group 611: 	370 
    -- CP-element group 611: 	378 
    -- CP-element group 611: 	382 
    -- CP-element group 611: 	390 
    -- CP-element group 611: 	401 
    -- CP-element group 611: 	405 
    -- CP-element group 611: 	409 
    -- CP-element group 611: 	417 
    -- CP-element group 611: 	421 
    -- CP-element group 611: 	429 
    -- CP-element group 611: 	449 
    -- CP-element group 611: 	465 
    -- CP-element group 611: 	473 
    -- CP-element group 611: 	477 
    -- CP-element group 611: 	481 
    -- CP-element group 611: 	485 
    -- CP-element group 611: 	493 
    -- CP-element group 611: 	497 
    -- CP-element group 611: 	501 
    -- CP-element group 611: 	505 
    -- CP-element group 611: 	509 
    -- CP-element group 611: 	513 
    -- CP-element group 611: 	517 
    -- CP-element group 611: 	521 
    -- CP-element group 611: 	525 
    -- CP-element group 611: 	529 
    -- CP-element group 611: 	533 
    -- CP-element group 611: 	537 
    -- CP-element group 611: 	541 
    -- CP-element group 611: 	549 
    -- CP-element group 611: 	553 
    -- CP-element group 611: 	557 
    -- CP-element group 611: 	561 
    -- CP-element group 611: 	565 
    -- CP-element group 611: 	571 
    -- CP-element group 611: 	572 
    -- CP-element group 611: 	576 
    -- CP-element group 611: 	580 
    -- CP-element group 611: 	600 
    -- CP-element group 611: successors 
    -- CP-element group 611: 	109 
    -- CP-element group 611:  members (1) 
      -- CP-element group 611: 	 branch_block_stmt_43/do_while_stmt_588/do_while_stmt_588_loop_body/$exit
      -- 
    zeropad_cp_element_group_611: block -- 
      constant place_capacities: IntegerArray(0 to 40) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15,16 => 15,17 => 15,18 => 15,19 => 15,20 => 15,21 => 15,22 => 15,23 => 15,24 => 15,25 => 15,26 => 15,27 => 15,28 => 15,29 => 15,30 => 15,31 => 15,32 => 15,33 => 15,34 => 15,35 => 15,36 => 15,37 => 15,38 => 15,39 => 15,40 => 15);
      constant place_markings: IntegerArray(0 to 40)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0,28 => 0,29 => 0,30 => 0,31 => 0,32 => 0,33 => 0,34 => 0,35 => 0,36 => 0,37 => 0,38 => 0,39 => 0,40 => 0);
      constant place_delays: IntegerArray(0 to 40) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0,28 => 0,29 => 0,30 => 0,31 => 0,32 => 0,33 => 0,34 => 0,35 => 0,36 => 0,37 => 0,38 => 0,39 => 0,40 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_611"; 
      signal preds: BooleanArray(1 to 41); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(354) & zeropad_CP_182_elements(358) & zeropad_CP_182_elements(370) & zeropad_CP_182_elements(378) & zeropad_CP_182_elements(382) & zeropad_CP_182_elements(390) & zeropad_CP_182_elements(401) & zeropad_CP_182_elements(405) & zeropad_CP_182_elements(409) & zeropad_CP_182_elements(417) & zeropad_CP_182_elements(421) & zeropad_CP_182_elements(429) & zeropad_CP_182_elements(449) & zeropad_CP_182_elements(465) & zeropad_CP_182_elements(473) & zeropad_CP_182_elements(477) & zeropad_CP_182_elements(481) & zeropad_CP_182_elements(485) & zeropad_CP_182_elements(493) & zeropad_CP_182_elements(497) & zeropad_CP_182_elements(501) & zeropad_CP_182_elements(505) & zeropad_CP_182_elements(509) & zeropad_CP_182_elements(513) & zeropad_CP_182_elements(517) & zeropad_CP_182_elements(521) & zeropad_CP_182_elements(525) & zeropad_CP_182_elements(529) & zeropad_CP_182_elements(533) & zeropad_CP_182_elements(537) & zeropad_CP_182_elements(541) & zeropad_CP_182_elements(549) & zeropad_CP_182_elements(553) & zeropad_CP_182_elements(557) & zeropad_CP_182_elements(561) & zeropad_CP_182_elements(565) & zeropad_CP_182_elements(571) & zeropad_CP_182_elements(572) & zeropad_CP_182_elements(576) & zeropad_CP_182_elements(580) & zeropad_CP_182_elements(600);
      gj_zeropad_cp_element_group_611 : generic_join generic map(name => joinName, number_of_predecessors => 41, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(611), clk => clk, reset => reset); --
    end block;
    -- CP-element group 612:  transition  input  bypass  pipeline-parent 
    -- CP-element group 612: predecessors 
    -- CP-element group 612: 	108 
    -- CP-element group 612: successors 
    -- CP-element group 612:  members (2) 
      -- CP-element group 612: 	 branch_block_stmt_43/do_while_stmt_588/loop_exit/$exit
      -- CP-element group 612: 	 branch_block_stmt_43/do_while_stmt_588/loop_exit/ack
      -- 
    ack_2607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 612_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_588_branch_ack_0, ack => zeropad_CP_182_elements(612)); -- 
    -- CP-element group 613:  transition  input  bypass  pipeline-parent 
    -- CP-element group 613: predecessors 
    -- CP-element group 613: 	108 
    -- CP-element group 613: successors 
    -- CP-element group 613:  members (2) 
      -- CP-element group 613: 	 branch_block_stmt_43/do_while_stmt_588/loop_taken/$exit
      -- CP-element group 613: 	 branch_block_stmt_43/do_while_stmt_588/loop_taken/ack
      -- 
    ack_2611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 613_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_588_branch_ack_1, ack => zeropad_CP_182_elements(613)); -- 
    -- CP-element group 614:  transition  bypass  pipeline-parent 
    -- CP-element group 614: predecessors 
    -- CP-element group 614: 	106 
    -- CP-element group 614: successors 
    -- CP-element group 614: 	1 
    -- CP-element group 614:  members (1) 
      -- CP-element group 614: 	 branch_block_stmt_43/do_while_stmt_588/$exit
      -- 
    zeropad_CP_182_elements(614) <= zeropad_CP_182_elements(106);
    -- CP-element group 615:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 615: predecessors 
    -- CP-element group 615: 	1 
    -- CP-element group 615: successors 
    -- CP-element group 615: 	617 
    -- CP-element group 615: 	618 
    -- CP-element group 615:  members (18) 
      -- CP-element group 615: 	 branch_block_stmt_43/merge_stmt_1336__exit__
      -- CP-element group 615: 	 branch_block_stmt_43/assign_stmt_1342__entry__
      -- CP-element group 615: 	 branch_block_stmt_43/if_stmt_1332_if_link/$exit
      -- CP-element group 615: 	 branch_block_stmt_43/if_stmt_1332_if_link/if_choice_transition
      -- CP-element group 615: 	 branch_block_stmt_43/ifx_xend253_whilex_xend
      -- CP-element group 615: 	 branch_block_stmt_43/assign_stmt_1342/$entry
      -- CP-element group 615: 	 branch_block_stmt_43/assign_stmt_1342/type_cast_1341_sample_start_
      -- CP-element group 615: 	 branch_block_stmt_43/assign_stmt_1342/type_cast_1341_update_start_
      -- CP-element group 615: 	 branch_block_stmt_43/assign_stmt_1342/type_cast_1341_Sample/$entry
      -- CP-element group 615: 	 branch_block_stmt_43/assign_stmt_1342/type_cast_1341_Sample/rr
      -- CP-element group 615: 	 branch_block_stmt_43/assign_stmt_1342/type_cast_1341_Update/$entry
      -- CP-element group 615: 	 branch_block_stmt_43/assign_stmt_1342/type_cast_1341_Update/cr
      -- CP-element group 615: 	 branch_block_stmt_43/ifx_xend253_whilex_xend_PhiReq/$entry
      -- CP-element group 615: 	 branch_block_stmt_43/ifx_xend253_whilex_xend_PhiReq/$exit
      -- CP-element group 615: 	 branch_block_stmt_43/merge_stmt_1336_PhiReqMerge
      -- CP-element group 615: 	 branch_block_stmt_43/merge_stmt_1336_PhiAck/$entry
      -- CP-element group 615: 	 branch_block_stmt_43/merge_stmt_1336_PhiAck/$exit
      -- CP-element group 615: 	 branch_block_stmt_43/merge_stmt_1336_PhiAck/dummy
      -- 
    if_choice_transition_2625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 615_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1332_branch_ack_1, ack => zeropad_CP_182_elements(615)); -- 
    rr_2641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(615), ack => type_cast_1341_inst_req_0); -- 
    cr_2646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(615), ack => type_cast_1341_inst_req_1); -- 
    -- CP-element group 616:  merge  transition  place  input  bypass 
    -- CP-element group 616: predecessors 
    -- CP-element group 616: 	1 
    -- CP-element group 616: successors 
    -- CP-element group 616:  members (5) 
      -- CP-element group 616: 	 branch_block_stmt_43/if_stmt_1332__exit__
      -- CP-element group 616: 	 branch_block_stmt_43/merge_stmt_1336__entry__
      -- CP-element group 616: 	 branch_block_stmt_43/if_stmt_1332_else_link/$exit
      -- CP-element group 616: 	 branch_block_stmt_43/if_stmt_1332_else_link/else_choice_transition
      -- CP-element group 616: 	 branch_block_stmt_43/merge_stmt_1336_dead_link/$entry
      -- 
    else_choice_transition_2629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 616_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1332_branch_ack_0, ack => zeropad_CP_182_elements(616)); -- 
    -- CP-element group 617:  transition  input  bypass 
    -- CP-element group 617: predecessors 
    -- CP-element group 617: 	615 
    -- CP-element group 617: successors 
    -- CP-element group 617:  members (3) 
      -- CP-element group 617: 	 branch_block_stmt_43/assign_stmt_1342/type_cast_1341_sample_completed_
      -- CP-element group 617: 	 branch_block_stmt_43/assign_stmt_1342/type_cast_1341_Sample/$exit
      -- CP-element group 617: 	 branch_block_stmt_43/assign_stmt_1342/type_cast_1341_Sample/ra
      -- 
    ra_2642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 617_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1341_inst_ack_0, ack => zeropad_CP_182_elements(617)); -- 
    -- CP-element group 618:  fork  transition  place  input  output  bypass 
    -- CP-element group 618: predecessors 
    -- CP-element group 618: 	615 
    -- CP-element group 618: successors 
    -- CP-element group 618: 	619 
    -- CP-element group 618: 	620 
    -- CP-element group 618: 	622 
    -- CP-element group 618: 	624 
    -- CP-element group 618: 	626 
    -- CP-element group 618: 	628 
    -- CP-element group 618: 	630 
    -- CP-element group 618: 	632 
    -- CP-element group 618: 	634 
    -- CP-element group 618: 	636 
    -- CP-element group 618: 	638 
    -- CP-element group 618:  members (40) 
      -- CP-element group 618: 	 branch_block_stmt_43/assign_stmt_1342__exit__
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453__entry__
      -- CP-element group 618: 	 branch_block_stmt_43/assign_stmt_1342/$exit
      -- CP-element group 618: 	 branch_block_stmt_43/assign_stmt_1342/type_cast_1341_update_completed_
      -- CP-element group 618: 	 branch_block_stmt_43/assign_stmt_1342/type_cast_1341_Update/$exit
      -- CP-element group 618: 	 branch_block_stmt_43/assign_stmt_1342/type_cast_1341_Update/ca
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/$entry
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/call_stmt_1345_sample_start_
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/call_stmt_1345_update_start_
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/call_stmt_1345_Sample/$entry
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/call_stmt_1345_Sample/crr
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/call_stmt_1345_Update/$entry
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/call_stmt_1345_Update/ccr
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1349_update_start_
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1349_Update/$entry
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1349_Update/cr
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1358_update_start_
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1358_Update/$entry
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1358_Update/cr
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1368_update_start_
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1368_Update/$entry
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1368_Update/cr
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1378_update_start_
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1378_Update/$entry
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1378_Update/cr
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1388_update_start_
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1388_Update/$entry
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1388_Update/cr
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1398_update_start_
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1398_Update/$entry
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1398_Update/cr
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1408_update_start_
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1408_Update/$entry
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1408_Update/cr
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1418_update_start_
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1418_Update/$entry
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1418_Update/cr
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1428_update_start_
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1428_Update/$entry
      -- CP-element group 618: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1428_Update/cr
      -- 
    ca_2647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 618_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1341_inst_ack_1, ack => zeropad_CP_182_elements(618)); -- 
    crr_2658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(618), ack => call_stmt_1345_call_req_0); -- 
    ccr_2663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(618), ack => call_stmt_1345_call_req_1); -- 
    cr_2677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(618), ack => type_cast_1349_inst_req_1); -- 
    cr_2691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(618), ack => type_cast_1358_inst_req_1); -- 
    cr_2705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(618), ack => type_cast_1368_inst_req_1); -- 
    cr_2719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(618), ack => type_cast_1378_inst_req_1); -- 
    cr_2733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(618), ack => type_cast_1388_inst_req_1); -- 
    cr_2747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(618), ack => type_cast_1398_inst_req_1); -- 
    cr_2761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(618), ack => type_cast_1408_inst_req_1); -- 
    cr_2775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(618), ack => type_cast_1418_inst_req_1); -- 
    cr_2789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(618), ack => type_cast_1428_inst_req_1); -- 
    -- CP-element group 619:  transition  input  bypass 
    -- CP-element group 619: predecessors 
    -- CP-element group 619: 	618 
    -- CP-element group 619: successors 
    -- CP-element group 619:  members (3) 
      -- CP-element group 619: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/call_stmt_1345_sample_completed_
      -- CP-element group 619: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/call_stmt_1345_Sample/$exit
      -- CP-element group 619: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/call_stmt_1345_Sample/cra
      -- 
    cra_2659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 619_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1345_call_ack_0, ack => zeropad_CP_182_elements(619)); -- 
    -- CP-element group 620:  transition  input  output  bypass 
    -- CP-element group 620: predecessors 
    -- CP-element group 620: 	618 
    -- CP-element group 620: successors 
    -- CP-element group 620: 	621 
    -- CP-element group 620:  members (6) 
      -- CP-element group 620: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/call_stmt_1345_update_completed_
      -- CP-element group 620: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/call_stmt_1345_Update/$exit
      -- CP-element group 620: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/call_stmt_1345_Update/cca
      -- CP-element group 620: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1349_sample_start_
      -- CP-element group 620: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1349_Sample/$entry
      -- CP-element group 620: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1349_Sample/rr
      -- 
    cca_2664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 620_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1345_call_ack_1, ack => zeropad_CP_182_elements(620)); -- 
    rr_2672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(620), ack => type_cast_1349_inst_req_0); -- 
    -- CP-element group 621:  transition  input  bypass 
    -- CP-element group 621: predecessors 
    -- CP-element group 621: 	620 
    -- CP-element group 621: successors 
    -- CP-element group 621:  members (3) 
      -- CP-element group 621: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1349_sample_completed_
      -- CP-element group 621: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1349_Sample/$exit
      -- CP-element group 621: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1349_Sample/ra
      -- 
    ra_2673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 621_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1349_inst_ack_0, ack => zeropad_CP_182_elements(621)); -- 
    -- CP-element group 622:  fork  transition  input  output  bypass 
    -- CP-element group 622: predecessors 
    -- CP-element group 622: 	618 
    -- CP-element group 622: successors 
    -- CP-element group 622: 	623 
    -- CP-element group 622: 	625 
    -- CP-element group 622: 	627 
    -- CP-element group 622: 	629 
    -- CP-element group 622: 	631 
    -- CP-element group 622: 	633 
    -- CP-element group 622: 	635 
    -- CP-element group 622: 	637 
    -- CP-element group 622:  members (27) 
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1349_update_completed_
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1349_Update/$exit
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1349_Update/ca
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1358_sample_start_
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1358_Sample/$entry
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1358_Sample/rr
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1368_sample_start_
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1368_Sample/$entry
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1368_Sample/rr
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1378_sample_start_
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1378_Sample/$entry
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1378_Sample/rr
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1388_sample_start_
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1388_Sample/$entry
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1388_Sample/rr
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1398_sample_start_
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1398_Sample/$entry
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1398_Sample/rr
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1408_sample_start_
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1408_Sample/$entry
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1408_Sample/rr
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1418_sample_start_
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1418_Sample/$entry
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1418_Sample/rr
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1428_sample_start_
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1428_Sample/$entry
      -- CP-element group 622: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1428_Sample/rr
      -- 
    ca_2678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 622_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1349_inst_ack_1, ack => zeropad_CP_182_elements(622)); -- 
    rr_2686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(622), ack => type_cast_1358_inst_req_0); -- 
    rr_2700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(622), ack => type_cast_1368_inst_req_0); -- 
    rr_2714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(622), ack => type_cast_1378_inst_req_0); -- 
    rr_2728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(622), ack => type_cast_1388_inst_req_0); -- 
    rr_2742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(622), ack => type_cast_1398_inst_req_0); -- 
    rr_2756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(622), ack => type_cast_1408_inst_req_0); -- 
    rr_2770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(622), ack => type_cast_1418_inst_req_0); -- 
    rr_2784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(622), ack => type_cast_1428_inst_req_0); -- 
    -- CP-element group 623:  transition  input  bypass 
    -- CP-element group 623: predecessors 
    -- CP-element group 623: 	622 
    -- CP-element group 623: successors 
    -- CP-element group 623:  members (3) 
      -- CP-element group 623: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1358_sample_completed_
      -- CP-element group 623: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1358_Sample/$exit
      -- CP-element group 623: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1358_Sample/ra
      -- 
    ra_2687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 623_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1358_inst_ack_0, ack => zeropad_CP_182_elements(623)); -- 
    -- CP-element group 624:  transition  input  bypass 
    -- CP-element group 624: predecessors 
    -- CP-element group 624: 	618 
    -- CP-element group 624: successors 
    -- CP-element group 624: 	659 
    -- CP-element group 624:  members (3) 
      -- CP-element group 624: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1358_update_completed_
      -- CP-element group 624: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1358_Update/$exit
      -- CP-element group 624: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1358_Update/ca
      -- 
    ca_2692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 624_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1358_inst_ack_1, ack => zeropad_CP_182_elements(624)); -- 
    -- CP-element group 625:  transition  input  bypass 
    -- CP-element group 625: predecessors 
    -- CP-element group 625: 	622 
    -- CP-element group 625: successors 
    -- CP-element group 625:  members (3) 
      -- CP-element group 625: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1368_sample_completed_
      -- CP-element group 625: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1368_Sample/$exit
      -- CP-element group 625: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1368_Sample/ra
      -- 
    ra_2701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 625_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1368_inst_ack_0, ack => zeropad_CP_182_elements(625)); -- 
    -- CP-element group 626:  transition  input  bypass 
    -- CP-element group 626: predecessors 
    -- CP-element group 626: 	618 
    -- CP-element group 626: successors 
    -- CP-element group 626: 	656 
    -- CP-element group 626:  members (3) 
      -- CP-element group 626: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1368_update_completed_
      -- CP-element group 626: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1368_Update/$exit
      -- CP-element group 626: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1368_Update/ca
      -- 
    ca_2706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 626_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1368_inst_ack_1, ack => zeropad_CP_182_elements(626)); -- 
    -- CP-element group 627:  transition  input  bypass 
    -- CP-element group 627: predecessors 
    -- CP-element group 627: 	622 
    -- CP-element group 627: successors 
    -- CP-element group 627:  members (3) 
      -- CP-element group 627: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1378_sample_completed_
      -- CP-element group 627: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1378_Sample/$exit
      -- CP-element group 627: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1378_Sample/ra
      -- 
    ra_2715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 627_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1378_inst_ack_0, ack => zeropad_CP_182_elements(627)); -- 
    -- CP-element group 628:  transition  input  bypass 
    -- CP-element group 628: predecessors 
    -- CP-element group 628: 	618 
    -- CP-element group 628: successors 
    -- CP-element group 628: 	653 
    -- CP-element group 628:  members (3) 
      -- CP-element group 628: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1378_update_completed_
      -- CP-element group 628: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1378_Update/$exit
      -- CP-element group 628: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1378_Update/ca
      -- 
    ca_2720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 628_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1378_inst_ack_1, ack => zeropad_CP_182_elements(628)); -- 
    -- CP-element group 629:  transition  input  bypass 
    -- CP-element group 629: predecessors 
    -- CP-element group 629: 	622 
    -- CP-element group 629: successors 
    -- CP-element group 629:  members (3) 
      -- CP-element group 629: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1388_sample_completed_
      -- CP-element group 629: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1388_Sample/$exit
      -- CP-element group 629: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1388_Sample/ra
      -- 
    ra_2729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 629_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1388_inst_ack_0, ack => zeropad_CP_182_elements(629)); -- 
    -- CP-element group 630:  transition  input  bypass 
    -- CP-element group 630: predecessors 
    -- CP-element group 630: 	618 
    -- CP-element group 630: successors 
    -- CP-element group 630: 	650 
    -- CP-element group 630:  members (3) 
      -- CP-element group 630: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1388_update_completed_
      -- CP-element group 630: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1388_Update/$exit
      -- CP-element group 630: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1388_Update/ca
      -- 
    ca_2734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 630_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1388_inst_ack_1, ack => zeropad_CP_182_elements(630)); -- 
    -- CP-element group 631:  transition  input  bypass 
    -- CP-element group 631: predecessors 
    -- CP-element group 631: 	622 
    -- CP-element group 631: successors 
    -- CP-element group 631:  members (3) 
      -- CP-element group 631: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1398_sample_completed_
      -- CP-element group 631: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1398_Sample/$exit
      -- CP-element group 631: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1398_Sample/ra
      -- 
    ra_2743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 631_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1398_inst_ack_0, ack => zeropad_CP_182_elements(631)); -- 
    -- CP-element group 632:  transition  input  bypass 
    -- CP-element group 632: predecessors 
    -- CP-element group 632: 	618 
    -- CP-element group 632: successors 
    -- CP-element group 632: 	647 
    -- CP-element group 632:  members (3) 
      -- CP-element group 632: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1398_update_completed_
      -- CP-element group 632: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1398_Update/$exit
      -- CP-element group 632: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1398_Update/ca
      -- 
    ca_2748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 632_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1398_inst_ack_1, ack => zeropad_CP_182_elements(632)); -- 
    -- CP-element group 633:  transition  input  bypass 
    -- CP-element group 633: predecessors 
    -- CP-element group 633: 	622 
    -- CP-element group 633: successors 
    -- CP-element group 633:  members (3) 
      -- CP-element group 633: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1408_sample_completed_
      -- CP-element group 633: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1408_Sample/$exit
      -- CP-element group 633: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1408_Sample/ra
      -- 
    ra_2757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 633_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1408_inst_ack_0, ack => zeropad_CP_182_elements(633)); -- 
    -- CP-element group 634:  transition  input  bypass 
    -- CP-element group 634: predecessors 
    -- CP-element group 634: 	618 
    -- CP-element group 634: successors 
    -- CP-element group 634: 	644 
    -- CP-element group 634:  members (3) 
      -- CP-element group 634: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1408_update_completed_
      -- CP-element group 634: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1408_Update/$exit
      -- CP-element group 634: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1408_Update/ca
      -- 
    ca_2762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 634_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1408_inst_ack_1, ack => zeropad_CP_182_elements(634)); -- 
    -- CP-element group 635:  transition  input  bypass 
    -- CP-element group 635: predecessors 
    -- CP-element group 635: 	622 
    -- CP-element group 635: successors 
    -- CP-element group 635:  members (3) 
      -- CP-element group 635: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1418_sample_completed_
      -- CP-element group 635: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1418_Sample/$exit
      -- CP-element group 635: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1418_Sample/ra
      -- 
    ra_2771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 635_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1418_inst_ack_0, ack => zeropad_CP_182_elements(635)); -- 
    -- CP-element group 636:  transition  input  bypass 
    -- CP-element group 636: predecessors 
    -- CP-element group 636: 	618 
    -- CP-element group 636: successors 
    -- CP-element group 636: 	641 
    -- CP-element group 636:  members (3) 
      -- CP-element group 636: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1418_update_completed_
      -- CP-element group 636: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1418_Update/$exit
      -- CP-element group 636: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1418_Update/ca
      -- 
    ca_2776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 636_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1418_inst_ack_1, ack => zeropad_CP_182_elements(636)); -- 
    -- CP-element group 637:  transition  input  bypass 
    -- CP-element group 637: predecessors 
    -- CP-element group 637: 	622 
    -- CP-element group 637: successors 
    -- CP-element group 637:  members (3) 
      -- CP-element group 637: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1428_sample_completed_
      -- CP-element group 637: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1428_Sample/$exit
      -- CP-element group 637: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1428_Sample/ra
      -- 
    ra_2785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 637_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1428_inst_ack_0, ack => zeropad_CP_182_elements(637)); -- 
    -- CP-element group 638:  transition  input  output  bypass 
    -- CP-element group 638: predecessors 
    -- CP-element group 638: 	618 
    -- CP-element group 638: successors 
    -- CP-element group 638: 	639 
    -- CP-element group 638:  members (6) 
      -- CP-element group 638: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1428_update_completed_
      -- CP-element group 638: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1428_Update/$exit
      -- CP-element group 638: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/type_cast_1428_Update/ca
      -- CP-element group 638: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1430_sample_start_
      -- CP-element group 638: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1430_Sample/$entry
      -- CP-element group 638: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1430_Sample/req
      -- 
    ca_2790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 638_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1428_inst_ack_1, ack => zeropad_CP_182_elements(638)); -- 
    req_2798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(638), ack => WPIPE_Zeropad_output_pipe_1430_inst_req_0); -- 
    -- CP-element group 639:  transition  input  output  bypass 
    -- CP-element group 639: predecessors 
    -- CP-element group 639: 	638 
    -- CP-element group 639: successors 
    -- CP-element group 639: 	640 
    -- CP-element group 639:  members (6) 
      -- CP-element group 639: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1430_Update/req
      -- CP-element group 639: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1430_Update/$entry
      -- CP-element group 639: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1430_sample_completed_
      -- CP-element group 639: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1430_update_start_
      -- CP-element group 639: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1430_Sample/$exit
      -- CP-element group 639: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1430_Sample/ack
      -- 
    ack_2799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 639_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1430_inst_ack_0, ack => zeropad_CP_182_elements(639)); -- 
    req_2803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(639), ack => WPIPE_Zeropad_output_pipe_1430_inst_req_1); -- 
    -- CP-element group 640:  transition  input  bypass 
    -- CP-element group 640: predecessors 
    -- CP-element group 640: 	639 
    -- CP-element group 640: successors 
    -- CP-element group 640: 	641 
    -- CP-element group 640:  members (3) 
      -- CP-element group 640: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1430_Update/ack
      -- CP-element group 640: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1430_Update/$exit
      -- CP-element group 640: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1430_update_completed_
      -- 
    ack_2804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 640_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1430_inst_ack_1, ack => zeropad_CP_182_elements(640)); -- 
    -- CP-element group 641:  join  transition  output  bypass 
    -- CP-element group 641: predecessors 
    -- CP-element group 641: 	636 
    -- CP-element group 641: 	640 
    -- CP-element group 641: successors 
    -- CP-element group 641: 	642 
    -- CP-element group 641:  members (3) 
      -- CP-element group 641: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1433_sample_start_
      -- CP-element group 641: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1433_Sample/$entry
      -- CP-element group 641: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1433_Sample/req
      -- 
    req_2812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(641), ack => WPIPE_Zeropad_output_pipe_1433_inst_req_0); -- 
    zeropad_cp_element_group_641: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_641"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(636) & zeropad_CP_182_elements(640);
      gj_zeropad_cp_element_group_641 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(641), clk => clk, reset => reset); --
    end block;
    -- CP-element group 642:  transition  input  output  bypass 
    -- CP-element group 642: predecessors 
    -- CP-element group 642: 	641 
    -- CP-element group 642: successors 
    -- CP-element group 642: 	643 
    -- CP-element group 642:  members (6) 
      -- CP-element group 642: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1433_update_start_
      -- CP-element group 642: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1433_sample_completed_
      -- CP-element group 642: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1433_Sample/$exit
      -- CP-element group 642: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1433_Sample/ack
      -- CP-element group 642: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1433_Update/$entry
      -- CP-element group 642: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1433_Update/req
      -- 
    ack_2813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 642_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1433_inst_ack_0, ack => zeropad_CP_182_elements(642)); -- 
    req_2817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(642), ack => WPIPE_Zeropad_output_pipe_1433_inst_req_1); -- 
    -- CP-element group 643:  transition  input  bypass 
    -- CP-element group 643: predecessors 
    -- CP-element group 643: 	642 
    -- CP-element group 643: successors 
    -- CP-element group 643: 	644 
    -- CP-element group 643:  members (3) 
      -- CP-element group 643: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1433_update_completed_
      -- CP-element group 643: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1433_Update/$exit
      -- CP-element group 643: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1433_Update/ack
      -- 
    ack_2818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 643_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1433_inst_ack_1, ack => zeropad_CP_182_elements(643)); -- 
    -- CP-element group 644:  join  transition  output  bypass 
    -- CP-element group 644: predecessors 
    -- CP-element group 644: 	634 
    -- CP-element group 644: 	643 
    -- CP-element group 644: successors 
    -- CP-element group 644: 	645 
    -- CP-element group 644:  members (3) 
      -- CP-element group 644: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1436_sample_start_
      -- CP-element group 644: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1436_Sample/$entry
      -- CP-element group 644: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1436_Sample/req
      -- 
    req_2826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(644), ack => WPIPE_Zeropad_output_pipe_1436_inst_req_0); -- 
    zeropad_cp_element_group_644: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_644"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(634) & zeropad_CP_182_elements(643);
      gj_zeropad_cp_element_group_644 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(644), clk => clk, reset => reset); --
    end block;
    -- CP-element group 645:  transition  input  output  bypass 
    -- CP-element group 645: predecessors 
    -- CP-element group 645: 	644 
    -- CP-element group 645: successors 
    -- CP-element group 645: 	646 
    -- CP-element group 645:  members (6) 
      -- CP-element group 645: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1436_Update/req
      -- CP-element group 645: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1436_sample_completed_
      -- CP-element group 645: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1436_update_start_
      -- CP-element group 645: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1436_Update/$entry
      -- CP-element group 645: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1436_Sample/ack
      -- CP-element group 645: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1436_Sample/$exit
      -- 
    ack_2827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 645_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1436_inst_ack_0, ack => zeropad_CP_182_elements(645)); -- 
    req_2831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(645), ack => WPIPE_Zeropad_output_pipe_1436_inst_req_1); -- 
    -- CP-element group 646:  transition  input  bypass 
    -- CP-element group 646: predecessors 
    -- CP-element group 646: 	645 
    -- CP-element group 646: successors 
    -- CP-element group 646: 	647 
    -- CP-element group 646:  members (3) 
      -- CP-element group 646: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1436_Update/ack
      -- CP-element group 646: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1436_update_completed_
      -- CP-element group 646: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1436_Update/$exit
      -- 
    ack_2832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 646_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1436_inst_ack_1, ack => zeropad_CP_182_elements(646)); -- 
    -- CP-element group 647:  join  transition  output  bypass 
    -- CP-element group 647: predecessors 
    -- CP-element group 647: 	632 
    -- CP-element group 647: 	646 
    -- CP-element group 647: successors 
    -- CP-element group 647: 	648 
    -- CP-element group 647:  members (3) 
      -- CP-element group 647: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1439_sample_start_
      -- CP-element group 647: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1439_Sample/$entry
      -- CP-element group 647: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1439_Sample/req
      -- 
    req_2840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(647), ack => WPIPE_Zeropad_output_pipe_1439_inst_req_0); -- 
    zeropad_cp_element_group_647: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_647"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(632) & zeropad_CP_182_elements(646);
      gj_zeropad_cp_element_group_647 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(647), clk => clk, reset => reset); --
    end block;
    -- CP-element group 648:  transition  input  output  bypass 
    -- CP-element group 648: predecessors 
    -- CP-element group 648: 	647 
    -- CP-element group 648: successors 
    -- CP-element group 648: 	649 
    -- CP-element group 648:  members (6) 
      -- CP-element group 648: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1439_sample_completed_
      -- CP-element group 648: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1439_update_start_
      -- CP-element group 648: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1439_Sample/$exit
      -- CP-element group 648: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1439_Sample/ack
      -- CP-element group 648: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1439_Update/req
      -- CP-element group 648: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1439_Update/$entry
      -- 
    ack_2841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 648_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1439_inst_ack_0, ack => zeropad_CP_182_elements(648)); -- 
    req_2845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(648), ack => WPIPE_Zeropad_output_pipe_1439_inst_req_1); -- 
    -- CP-element group 649:  transition  input  bypass 
    -- CP-element group 649: predecessors 
    -- CP-element group 649: 	648 
    -- CP-element group 649: successors 
    -- CP-element group 649: 	650 
    -- CP-element group 649:  members (3) 
      -- CP-element group 649: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1439_update_completed_
      -- CP-element group 649: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1439_Update/ack
      -- CP-element group 649: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1439_Update/$exit
      -- 
    ack_2846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 649_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1439_inst_ack_1, ack => zeropad_CP_182_elements(649)); -- 
    -- CP-element group 650:  join  transition  output  bypass 
    -- CP-element group 650: predecessors 
    -- CP-element group 650: 	630 
    -- CP-element group 650: 	649 
    -- CP-element group 650: successors 
    -- CP-element group 650: 	651 
    -- CP-element group 650:  members (3) 
      -- CP-element group 650: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1442_Sample/$entry
      -- CP-element group 650: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1442_Sample/req
      -- CP-element group 650: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1442_sample_start_
      -- 
    req_2854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(650), ack => WPIPE_Zeropad_output_pipe_1442_inst_req_0); -- 
    zeropad_cp_element_group_650: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_650"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(630) & zeropad_CP_182_elements(649);
      gj_zeropad_cp_element_group_650 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(650), clk => clk, reset => reset); --
    end block;
    -- CP-element group 651:  transition  input  output  bypass 
    -- CP-element group 651: predecessors 
    -- CP-element group 651: 	650 
    -- CP-element group 651: successors 
    -- CP-element group 651: 	652 
    -- CP-element group 651:  members (6) 
      -- CP-element group 651: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1442_sample_completed_
      -- CP-element group 651: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1442_Sample/$exit
      -- CP-element group 651: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1442_update_start_
      -- CP-element group 651: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1442_Sample/ack
      -- CP-element group 651: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1442_Update/$entry
      -- CP-element group 651: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1442_Update/req
      -- 
    ack_2855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 651_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1442_inst_ack_0, ack => zeropad_CP_182_elements(651)); -- 
    req_2859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(651), ack => WPIPE_Zeropad_output_pipe_1442_inst_req_1); -- 
    -- CP-element group 652:  transition  input  bypass 
    -- CP-element group 652: predecessors 
    -- CP-element group 652: 	651 
    -- CP-element group 652: successors 
    -- CP-element group 652: 	653 
    -- CP-element group 652:  members (3) 
      -- CP-element group 652: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1442_update_completed_
      -- CP-element group 652: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1442_Update/$exit
      -- CP-element group 652: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1442_Update/ack
      -- 
    ack_2860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 652_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1442_inst_ack_1, ack => zeropad_CP_182_elements(652)); -- 
    -- CP-element group 653:  join  transition  output  bypass 
    -- CP-element group 653: predecessors 
    -- CP-element group 653: 	628 
    -- CP-element group 653: 	652 
    -- CP-element group 653: successors 
    -- CP-element group 653: 	654 
    -- CP-element group 653:  members (3) 
      -- CP-element group 653: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1445_Sample/req
      -- CP-element group 653: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1445_sample_start_
      -- CP-element group 653: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1445_Sample/$entry
      -- 
    req_2868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(653), ack => WPIPE_Zeropad_output_pipe_1445_inst_req_0); -- 
    zeropad_cp_element_group_653: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_653"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(628) & zeropad_CP_182_elements(652);
      gj_zeropad_cp_element_group_653 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(653), clk => clk, reset => reset); --
    end block;
    -- CP-element group 654:  transition  input  output  bypass 
    -- CP-element group 654: predecessors 
    -- CP-element group 654: 	653 
    -- CP-element group 654: successors 
    -- CP-element group 654: 	655 
    -- CP-element group 654:  members (6) 
      -- CP-element group 654: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1445_Sample/$exit
      -- CP-element group 654: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1445_Sample/ack
      -- CP-element group 654: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1445_Update/$entry
      -- CP-element group 654: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1445_Update/req
      -- CP-element group 654: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1445_sample_completed_
      -- CP-element group 654: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1445_update_start_
      -- 
    ack_2869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 654_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1445_inst_ack_0, ack => zeropad_CP_182_elements(654)); -- 
    req_2873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(654), ack => WPIPE_Zeropad_output_pipe_1445_inst_req_1); -- 
    -- CP-element group 655:  transition  input  bypass 
    -- CP-element group 655: predecessors 
    -- CP-element group 655: 	654 
    -- CP-element group 655: successors 
    -- CP-element group 655: 	656 
    -- CP-element group 655:  members (3) 
      -- CP-element group 655: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1445_Update/$exit
      -- CP-element group 655: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1445_Update/ack
      -- CP-element group 655: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1445_update_completed_
      -- 
    ack_2874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 655_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1445_inst_ack_1, ack => zeropad_CP_182_elements(655)); -- 
    -- CP-element group 656:  join  transition  output  bypass 
    -- CP-element group 656: predecessors 
    -- CP-element group 656: 	626 
    -- CP-element group 656: 	655 
    -- CP-element group 656: successors 
    -- CP-element group 656: 	657 
    -- CP-element group 656:  members (3) 
      -- CP-element group 656: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1448_sample_start_
      -- CP-element group 656: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1448_Sample/$entry
      -- CP-element group 656: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1448_Sample/req
      -- 
    req_2882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(656), ack => WPIPE_Zeropad_output_pipe_1448_inst_req_0); -- 
    zeropad_cp_element_group_656: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_656"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(626) & zeropad_CP_182_elements(655);
      gj_zeropad_cp_element_group_656 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(656), clk => clk, reset => reset); --
    end block;
    -- CP-element group 657:  transition  input  output  bypass 
    -- CP-element group 657: predecessors 
    -- CP-element group 657: 	656 
    -- CP-element group 657: successors 
    -- CP-element group 657: 	658 
    -- CP-element group 657:  members (6) 
      -- CP-element group 657: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1448_sample_completed_
      -- CP-element group 657: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1448_update_start_
      -- CP-element group 657: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1448_Sample/$exit
      -- CP-element group 657: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1448_Update/req
      -- CP-element group 657: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1448_Update/$entry
      -- CP-element group 657: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1448_Sample/ack
      -- 
    ack_2883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 657_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1448_inst_ack_0, ack => zeropad_CP_182_elements(657)); -- 
    req_2887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(657), ack => WPIPE_Zeropad_output_pipe_1448_inst_req_1); -- 
    -- CP-element group 658:  transition  input  bypass 
    -- CP-element group 658: predecessors 
    -- CP-element group 658: 	657 
    -- CP-element group 658: successors 
    -- CP-element group 658: 	659 
    -- CP-element group 658:  members (3) 
      -- CP-element group 658: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1448_update_completed_
      -- CP-element group 658: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1448_Update/ack
      -- CP-element group 658: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1448_Update/$exit
      -- 
    ack_2888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 658_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1448_inst_ack_1, ack => zeropad_CP_182_elements(658)); -- 
    -- CP-element group 659:  join  transition  output  bypass 
    -- CP-element group 659: predecessors 
    -- CP-element group 659: 	624 
    -- CP-element group 659: 	658 
    -- CP-element group 659: successors 
    -- CP-element group 659: 	660 
    -- CP-element group 659:  members (3) 
      -- CP-element group 659: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1451_Sample/req
      -- CP-element group 659: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1451_Sample/$entry
      -- CP-element group 659: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1451_sample_start_
      -- 
    req_2896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(659), ack => WPIPE_Zeropad_output_pipe_1451_inst_req_0); -- 
    zeropad_cp_element_group_659: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_659"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(624) & zeropad_CP_182_elements(658);
      gj_zeropad_cp_element_group_659 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(659), clk => clk, reset => reset); --
    end block;
    -- CP-element group 660:  transition  input  output  bypass 
    -- CP-element group 660: predecessors 
    -- CP-element group 660: 	659 
    -- CP-element group 660: successors 
    -- CP-element group 660: 	661 
    -- CP-element group 660:  members (6) 
      -- CP-element group 660: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1451_Sample/ack
      -- CP-element group 660: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1451_Update/$entry
      -- CP-element group 660: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1451_Update/req
      -- CP-element group 660: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1451_Sample/$exit
      -- CP-element group 660: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1451_update_start_
      -- CP-element group 660: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1451_sample_completed_
      -- 
    ack_2897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 660_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1451_inst_ack_0, ack => zeropad_CP_182_elements(660)); -- 
    req_2901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(660), ack => WPIPE_Zeropad_output_pipe_1451_inst_req_1); -- 
    -- CP-element group 661:  branch  transition  place  input  output  bypass 
    -- CP-element group 661: predecessors 
    -- CP-element group 661: 	660 
    -- CP-element group 661: successors 
    -- CP-element group 661: 	662 
    -- CP-element group 661: 	663 
    -- CP-element group 661:  members (17) 
      -- CP-element group 661: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453__exit__
      -- CP-element group 661: 	 branch_block_stmt_43/assign_stmt_1460__entry__
      -- CP-element group 661: 	 branch_block_stmt_43/assign_stmt_1460__exit__
      -- CP-element group 661: 	 branch_block_stmt_43/if_stmt_1461__entry__
      -- CP-element group 661: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1451_Update/$exit
      -- CP-element group 661: 	 branch_block_stmt_43/assign_stmt_1460/$entry
      -- CP-element group 661: 	 branch_block_stmt_43/assign_stmt_1460/$exit
      -- CP-element group 661: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1451_Update/ack
      -- CP-element group 661: 	 branch_block_stmt_43/if_stmt_1461_dead_link/$entry
      -- CP-element group 661: 	 branch_block_stmt_43/if_stmt_1461_eval_test/$entry
      -- CP-element group 661: 	 branch_block_stmt_43/if_stmt_1461_eval_test/$exit
      -- CP-element group 661: 	 branch_block_stmt_43/if_stmt_1461_eval_test/branch_req
      -- CP-element group 661: 	 branch_block_stmt_43/if_stmt_1461_if_link/$entry
      -- CP-element group 661: 	 branch_block_stmt_43/if_stmt_1461_else_link/$entry
      -- CP-element group 661: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/WPIPE_Zeropad_output_pipe_1451_update_completed_
      -- CP-element group 661: 	 branch_block_stmt_43/call_stmt_1345_to_assign_stmt_1453/$exit
      -- CP-element group 661: 	 branch_block_stmt_43/R_cmp369459_1462_place
      -- 
    ack_2902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 661_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1451_inst_ack_1, ack => zeropad_CP_182_elements(661)); -- 
    branch_req_2913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(661), ack => if_stmt_1461_branch_req_0); -- 
    -- CP-element group 662:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 662: predecessors 
    -- CP-element group 662: 	661 
    -- CP-element group 662: successors 
    -- CP-element group 662: 	664 
    -- CP-element group 662: 	665 
    -- CP-element group 662: 	666 
    -- CP-element group 662: 	667 
    -- CP-element group 662:  members (24) 
      -- CP-element group 662: 	 branch_block_stmt_43/merge_stmt_1467__exit__
      -- CP-element group 662: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504__entry__
      -- CP-element group 662: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1470_Update/$entry
      -- CP-element group 662: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1470_Sample/rr
      -- CP-element group 662: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1470_Update/cr
      -- CP-element group 662: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1479_sample_start_
      -- CP-element group 662: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1479_update_start_
      -- CP-element group 662: 	 branch_block_stmt_43/if_stmt_1461_if_link/$exit
      -- CP-element group 662: 	 branch_block_stmt_43/if_stmt_1461_if_link/if_choice_transition
      -- CP-element group 662: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1470_Sample/$entry
      -- CP-element group 662: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1470_update_start_
      -- CP-element group 662: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1470_sample_start_
      -- CP-element group 662: 	 branch_block_stmt_43/whilex_xend_bbx_xnph
      -- CP-element group 662: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/$entry
      -- CP-element group 662: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1479_Update/cr
      -- CP-element group 662: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1479_Update/$entry
      -- CP-element group 662: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1479_Sample/rr
      -- CP-element group 662: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1479_Sample/$entry
      -- CP-element group 662: 	 branch_block_stmt_43/whilex_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 662: 	 branch_block_stmt_43/whilex_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 662: 	 branch_block_stmt_43/merge_stmt_1467_PhiReqMerge
      -- CP-element group 662: 	 branch_block_stmt_43/merge_stmt_1467_PhiAck/$entry
      -- CP-element group 662: 	 branch_block_stmt_43/merge_stmt_1467_PhiAck/$exit
      -- CP-element group 662: 	 branch_block_stmt_43/merge_stmt_1467_PhiAck/dummy
      -- 
    if_choice_transition_2918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 662_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1461_branch_ack_1, ack => zeropad_CP_182_elements(662)); -- 
    rr_2935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(662), ack => type_cast_1470_inst_req_0); -- 
    cr_2940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(662), ack => type_cast_1470_inst_req_1); -- 
    cr_2954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(662), ack => type_cast_1479_inst_req_1); -- 
    rr_2949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(662), ack => type_cast_1479_inst_req_0); -- 
    -- CP-element group 663:  transition  place  input  bypass 
    -- CP-element group 663: predecessors 
    -- CP-element group 663: 	661 
    -- CP-element group 663: successors 
    -- CP-element group 663: 	740 
    -- CP-element group 663:  members (5) 
      -- CP-element group 663: 	 branch_block_stmt_43/whilex_xend_forx_xend443
      -- CP-element group 663: 	 branch_block_stmt_43/if_stmt_1461_else_link/else_choice_transition
      -- CP-element group 663: 	 branch_block_stmt_43/if_stmt_1461_else_link/$exit
      -- CP-element group 663: 	 branch_block_stmt_43/whilex_xend_forx_xend443_PhiReq/$entry
      -- CP-element group 663: 	 branch_block_stmt_43/whilex_xend_forx_xend443_PhiReq/$exit
      -- 
    else_choice_transition_2922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 663_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1461_branch_ack_0, ack => zeropad_CP_182_elements(663)); -- 
    -- CP-element group 664:  transition  input  bypass 
    -- CP-element group 664: predecessors 
    -- CP-element group 664: 	662 
    -- CP-element group 664: successors 
    -- CP-element group 664:  members (3) 
      -- CP-element group 664: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1470_Sample/ra
      -- CP-element group 664: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1470_Sample/$exit
      -- CP-element group 664: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1470_sample_completed_
      -- 
    ra_2936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 664_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1470_inst_ack_0, ack => zeropad_CP_182_elements(664)); -- 
    -- CP-element group 665:  transition  input  bypass 
    -- CP-element group 665: predecessors 
    -- CP-element group 665: 	662 
    -- CP-element group 665: successors 
    -- CP-element group 665: 	668 
    -- CP-element group 665:  members (3) 
      -- CP-element group 665: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1470_Update/ca
      -- CP-element group 665: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1470_Update/$exit
      -- CP-element group 665: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1470_update_completed_
      -- 
    ca_2941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 665_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1470_inst_ack_1, ack => zeropad_CP_182_elements(665)); -- 
    -- CP-element group 666:  transition  input  bypass 
    -- CP-element group 666: predecessors 
    -- CP-element group 666: 	662 
    -- CP-element group 666: successors 
    -- CP-element group 666:  members (3) 
      -- CP-element group 666: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1479_sample_completed_
      -- CP-element group 666: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1479_Sample/ra
      -- CP-element group 666: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1479_Sample/$exit
      -- 
    ra_2950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 666_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1479_inst_ack_0, ack => zeropad_CP_182_elements(666)); -- 
    -- CP-element group 667:  transition  input  bypass 
    -- CP-element group 667: predecessors 
    -- CP-element group 667: 	662 
    -- CP-element group 667: successors 
    -- CP-element group 667: 	668 
    -- CP-element group 667:  members (3) 
      -- CP-element group 667: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1479_Update/ca
      -- CP-element group 667: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1479_Update/$exit
      -- CP-element group 667: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/type_cast_1479_update_completed_
      -- 
    ca_2955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 667_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1479_inst_ack_1, ack => zeropad_CP_182_elements(667)); -- 
    -- CP-element group 668:  join  transition  place  bypass 
    -- CP-element group 668: predecessors 
    -- CP-element group 668: 	665 
    -- CP-element group 668: 	667 
    -- CP-element group 668: successors 
    -- CP-element group 668: 	734 
    -- CP-element group 668:  members (6) 
      -- CP-element group 668: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504__exit__
      -- CP-element group 668: 	 branch_block_stmt_43/bbx_xnph_forx_xbody371
      -- CP-element group 668: 	 branch_block_stmt_43/assign_stmt_1471_to_assign_stmt_1504/$exit
      -- CP-element group 668: 	 branch_block_stmt_43/bbx_xnph_forx_xbody371_PhiReq/$entry
      -- CP-element group 668: 	 branch_block_stmt_43/bbx_xnph_forx_xbody371_PhiReq/phi_stmt_1507/$entry
      -- CP-element group 668: 	 branch_block_stmt_43/bbx_xnph_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/$entry
      -- 
    zeropad_cp_element_group_668: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_668"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(665) & zeropad_CP_182_elements(667);
      gj_zeropad_cp_element_group_668 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(668), clk => clk, reset => reset); --
    end block;
    -- CP-element group 669:  transition  input  bypass 
    -- CP-element group 669: predecessors 
    -- CP-element group 669: 	739 
    -- CP-element group 669: successors 
    -- CP-element group 669: 	714 
    -- CP-element group 669:  members (3) 
      -- CP-element group 669: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_final_index_sum_regn_sample_complete
      -- CP-element group 669: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_final_index_sum_regn_Sample/ack
      -- CP-element group 669: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_final_index_sum_regn_Sample/$exit
      -- 
    ack_2984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 669_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1521_index_offset_ack_0, ack => zeropad_CP_182_elements(669)); -- 
    -- CP-element group 670:  transition  input  output  bypass 
    -- CP-element group 670: predecessors 
    -- CP-element group 670: 	739 
    -- CP-element group 670: successors 
    -- CP-element group 670: 	671 
    -- CP-element group 670:  members (11) 
      -- CP-element group 670: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_final_index_sum_regn_Update/$exit
      -- CP-element group 670: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_final_index_sum_regn_Update/ack
      -- CP-element group 670: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_base_plus_offset/$entry
      -- CP-element group 670: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_base_plus_offset/$exit
      -- CP-element group 670: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_base_plus_offset/sum_rename_req
      -- CP-element group 670: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_base_plus_offset/sum_rename_ack
      -- CP-element group 670: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/addr_of_1522_request/$entry
      -- CP-element group 670: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/addr_of_1522_request/req
      -- CP-element group 670: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_offset_calculated
      -- CP-element group 670: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_root_address_calculated
      -- CP-element group 670: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/addr_of_1522_sample_start_
      -- 
    ack_2989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 670_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1521_index_offset_ack_1, ack => zeropad_CP_182_elements(670)); -- 
    req_2998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(670), ack => addr_of_1522_final_reg_req_0); -- 
    -- CP-element group 671:  transition  input  bypass 
    -- CP-element group 671: predecessors 
    -- CP-element group 671: 	670 
    -- CP-element group 671: successors 
    -- CP-element group 671:  members (3) 
      -- CP-element group 671: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/addr_of_1522_request/$exit
      -- CP-element group 671: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/addr_of_1522_request/ack
      -- CP-element group 671: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/addr_of_1522_sample_completed_
      -- 
    ack_2999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 671_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1522_final_reg_ack_0, ack => zeropad_CP_182_elements(671)); -- 
    -- CP-element group 672:  join  fork  transition  input  output  bypass 
    -- CP-element group 672: predecessors 
    -- CP-element group 672: 	739 
    -- CP-element group 672: successors 
    -- CP-element group 672: 	673 
    -- CP-element group 672:  members (24) 
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/addr_of_1522_complete/$exit
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/addr_of_1522_complete/ack
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_sample_start_
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Sample/word_access_start/word_0/rr
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Sample/word_access_start/word_0/$entry
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Sample/word_access_start/$entry
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Sample/$entry
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_word_addrgen/root_register_ack
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_word_addrgen/root_register_req
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_word_addrgen/$exit
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_word_addrgen/$entry
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/addr_of_1522_update_completed_
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_base_plus_offset/sum_rename_ack
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_base_plus_offset/sum_rename_req
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_base_plus_offset/$exit
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_base_plus_offset/$entry
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_base_addr_resize/base_resize_ack
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_base_addr_resize/base_resize_req
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_base_addr_resize/$exit
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_base_addr_resize/$entry
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_base_address_resized
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_root_address_calculated
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_word_address_calculated
      -- CP-element group 672: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_base_address_calculated
      -- 
    ack_3004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 672_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1522_final_reg_ack_1, ack => zeropad_CP_182_elements(672)); -- 
    rr_3037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(672), ack => ptr_deref_1526_load_0_req_0); -- 
    -- CP-element group 673:  transition  input  bypass 
    -- CP-element group 673: predecessors 
    -- CP-element group 673: 	672 
    -- CP-element group 673: successors 
    -- CP-element group 673:  members (5) 
      -- CP-element group 673: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_sample_completed_
      -- CP-element group 673: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Sample/word_access_start/word_0/ra
      -- CP-element group 673: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Sample/word_access_start/word_0/$exit
      -- CP-element group 673: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Sample/word_access_start/$exit
      -- CP-element group 673: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Sample/$exit
      -- 
    ra_3038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 673_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1526_load_0_ack_0, ack => zeropad_CP_182_elements(673)); -- 
    -- CP-element group 674:  fork  transition  input  output  bypass 
    -- CP-element group 674: predecessors 
    -- CP-element group 674: 	739 
    -- CP-element group 674: successors 
    -- CP-element group 674: 	675 
    -- CP-element group 674: 	677 
    -- CP-element group 674: 	679 
    -- CP-element group 674: 	681 
    -- CP-element group 674: 	683 
    -- CP-element group 674: 	685 
    -- CP-element group 674: 	687 
    -- CP-element group 674: 	689 
    -- CP-element group 674:  members (33) 
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1550_Sample/$entry
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1540_sample_start_
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Update/word_access_complete/word_0/$exit
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1590_sample_start_
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1550_sample_start_
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Update/word_access_complete/$exit
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_update_completed_
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Update/$exit
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1590_Sample/$entry
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1590_Sample/rr
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1550_Sample/rr
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Update/word_access_complete/word_0/ca
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1600_sample_start_
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Update/ptr_deref_1526_Merge/$entry
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Update/ptr_deref_1526_Merge/$exit
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1600_Sample/$entry
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Update/ptr_deref_1526_Merge/merge_req
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Update/ptr_deref_1526_Merge/merge_ack
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1530_sample_start_
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1600_Sample/rr
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1560_sample_start_
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1530_Sample/$entry
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1580_Sample/rr
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1580_sample_start_
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1570_Sample/rr
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1540_Sample/rr
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1570_Sample/$entry
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1570_sample_start_
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1540_Sample/$entry
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1580_Sample/$entry
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1530_Sample/rr
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1560_Sample/rr
      -- CP-element group 674: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1560_Sample/$entry
      -- 
    ca_3049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 674_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1526_load_0_ack_1, ack => zeropad_CP_182_elements(674)); -- 
    rr_3062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(674), ack => type_cast_1530_inst_req_0); -- 
    rr_3076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(674), ack => type_cast_1540_inst_req_0); -- 
    rr_3090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(674), ack => type_cast_1550_inst_req_0); -- 
    rr_3104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(674), ack => type_cast_1560_inst_req_0); -- 
    rr_3118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(674), ack => type_cast_1570_inst_req_0); -- 
    rr_3132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(674), ack => type_cast_1580_inst_req_0); -- 
    rr_3146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(674), ack => type_cast_1590_inst_req_0); -- 
    rr_3160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(674), ack => type_cast_1600_inst_req_0); -- 
    -- CP-element group 675:  transition  input  bypass 
    -- CP-element group 675: predecessors 
    -- CP-element group 675: 	674 
    -- CP-element group 675: successors 
    -- CP-element group 675:  members (3) 
      -- CP-element group 675: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1530_Sample/ra
      -- CP-element group 675: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1530_sample_completed_
      -- CP-element group 675: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1530_Sample/$exit
      -- 
    ra_3063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 675_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1530_inst_ack_0, ack => zeropad_CP_182_elements(675)); -- 
    -- CP-element group 676:  transition  input  bypass 
    -- CP-element group 676: predecessors 
    -- CP-element group 676: 	739 
    -- CP-element group 676: successors 
    -- CP-element group 676: 	711 
    -- CP-element group 676:  members (3) 
      -- CP-element group 676: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1530_Update/$exit
      -- CP-element group 676: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1530_Update/ca
      -- CP-element group 676: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1530_update_completed_
      -- 
    ca_3068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 676_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1530_inst_ack_1, ack => zeropad_CP_182_elements(676)); -- 
    -- CP-element group 677:  transition  input  bypass 
    -- CP-element group 677: predecessors 
    -- CP-element group 677: 	674 
    -- CP-element group 677: successors 
    -- CP-element group 677:  members (3) 
      -- CP-element group 677: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1540_sample_completed_
      -- CP-element group 677: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1540_Sample/ra
      -- CP-element group 677: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1540_Sample/$exit
      -- 
    ra_3077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 677_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1540_inst_ack_0, ack => zeropad_CP_182_elements(677)); -- 
    -- CP-element group 678:  transition  input  bypass 
    -- CP-element group 678: predecessors 
    -- CP-element group 678: 	739 
    -- CP-element group 678: successors 
    -- CP-element group 678: 	708 
    -- CP-element group 678:  members (3) 
      -- CP-element group 678: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1540_Update/ca
      -- CP-element group 678: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1540_Update/$exit
      -- CP-element group 678: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1540_update_completed_
      -- 
    ca_3082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 678_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1540_inst_ack_1, ack => zeropad_CP_182_elements(678)); -- 
    -- CP-element group 679:  transition  input  bypass 
    -- CP-element group 679: predecessors 
    -- CP-element group 679: 	674 
    -- CP-element group 679: successors 
    -- CP-element group 679:  members (3) 
      -- CP-element group 679: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1550_sample_completed_
      -- CP-element group 679: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1550_Sample/$exit
      -- CP-element group 679: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1550_Sample/ra
      -- 
    ra_3091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 679_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1550_inst_ack_0, ack => zeropad_CP_182_elements(679)); -- 
    -- CP-element group 680:  transition  input  bypass 
    -- CP-element group 680: predecessors 
    -- CP-element group 680: 	739 
    -- CP-element group 680: successors 
    -- CP-element group 680: 	705 
    -- CP-element group 680:  members (3) 
      -- CP-element group 680: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1550_update_completed_
      -- CP-element group 680: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1550_Update/$exit
      -- CP-element group 680: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1550_Update/ca
      -- 
    ca_3096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 680_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1550_inst_ack_1, ack => zeropad_CP_182_elements(680)); -- 
    -- CP-element group 681:  transition  input  bypass 
    -- CP-element group 681: predecessors 
    -- CP-element group 681: 	674 
    -- CP-element group 681: successors 
    -- CP-element group 681:  members (3) 
      -- CP-element group 681: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1560_sample_completed_
      -- CP-element group 681: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1560_Sample/ra
      -- CP-element group 681: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1560_Sample/$exit
      -- 
    ra_3105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 681_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1560_inst_ack_0, ack => zeropad_CP_182_elements(681)); -- 
    -- CP-element group 682:  transition  input  bypass 
    -- CP-element group 682: predecessors 
    -- CP-element group 682: 	739 
    -- CP-element group 682: successors 
    -- CP-element group 682: 	702 
    -- CP-element group 682:  members (3) 
      -- CP-element group 682: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1560_Update/ca
      -- CP-element group 682: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1560_Update/$exit
      -- CP-element group 682: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1560_update_completed_
      -- 
    ca_3110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 682_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1560_inst_ack_1, ack => zeropad_CP_182_elements(682)); -- 
    -- CP-element group 683:  transition  input  bypass 
    -- CP-element group 683: predecessors 
    -- CP-element group 683: 	674 
    -- CP-element group 683: successors 
    -- CP-element group 683:  members (3) 
      -- CP-element group 683: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1570_Sample/ra
      -- CP-element group 683: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1570_Sample/$exit
      -- CP-element group 683: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1570_sample_completed_
      -- 
    ra_3119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 683_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1570_inst_ack_0, ack => zeropad_CP_182_elements(683)); -- 
    -- CP-element group 684:  transition  input  bypass 
    -- CP-element group 684: predecessors 
    -- CP-element group 684: 	739 
    -- CP-element group 684: successors 
    -- CP-element group 684: 	699 
    -- CP-element group 684:  members (3) 
      -- CP-element group 684: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1570_Update/ca
      -- CP-element group 684: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1570_Update/$exit
      -- CP-element group 684: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1570_update_completed_
      -- 
    ca_3124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 684_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1570_inst_ack_1, ack => zeropad_CP_182_elements(684)); -- 
    -- CP-element group 685:  transition  input  bypass 
    -- CP-element group 685: predecessors 
    -- CP-element group 685: 	674 
    -- CP-element group 685: successors 
    -- CP-element group 685:  members (3) 
      -- CP-element group 685: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1580_Sample/ra
      -- CP-element group 685: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1580_Sample/$exit
      -- CP-element group 685: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1580_sample_completed_
      -- 
    ra_3133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 685_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1580_inst_ack_0, ack => zeropad_CP_182_elements(685)); -- 
    -- CP-element group 686:  transition  input  bypass 
    -- CP-element group 686: predecessors 
    -- CP-element group 686: 	739 
    -- CP-element group 686: successors 
    -- CP-element group 686: 	696 
    -- CP-element group 686:  members (3) 
      -- CP-element group 686: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1580_Update/ca
      -- CP-element group 686: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1580_Update/$exit
      -- CP-element group 686: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1580_update_completed_
      -- 
    ca_3138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 686_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1580_inst_ack_1, ack => zeropad_CP_182_elements(686)); -- 
    -- CP-element group 687:  transition  input  bypass 
    -- CP-element group 687: predecessors 
    -- CP-element group 687: 	674 
    -- CP-element group 687: successors 
    -- CP-element group 687:  members (3) 
      -- CP-element group 687: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1590_sample_completed_
      -- CP-element group 687: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1590_Sample/$exit
      -- CP-element group 687: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1590_Sample/ra
      -- 
    ra_3147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 687_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1590_inst_ack_0, ack => zeropad_CP_182_elements(687)); -- 
    -- CP-element group 688:  transition  input  bypass 
    -- CP-element group 688: predecessors 
    -- CP-element group 688: 	739 
    -- CP-element group 688: successors 
    -- CP-element group 688: 	693 
    -- CP-element group 688:  members (3) 
      -- CP-element group 688: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1590_update_completed_
      -- CP-element group 688: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1590_Update/ca
      -- CP-element group 688: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1590_Update/$exit
      -- 
    ca_3152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 688_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1590_inst_ack_1, ack => zeropad_CP_182_elements(688)); -- 
    -- CP-element group 689:  transition  input  bypass 
    -- CP-element group 689: predecessors 
    -- CP-element group 689: 	674 
    -- CP-element group 689: successors 
    -- CP-element group 689:  members (3) 
      -- CP-element group 689: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1600_sample_completed_
      -- CP-element group 689: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1600_Sample/$exit
      -- CP-element group 689: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1600_Sample/ra
      -- 
    ra_3161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 689_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1600_inst_ack_0, ack => zeropad_CP_182_elements(689)); -- 
    -- CP-element group 690:  transition  input  output  bypass 
    -- CP-element group 690: predecessors 
    -- CP-element group 690: 	739 
    -- CP-element group 690: successors 
    -- CP-element group 690: 	691 
    -- CP-element group 690:  members (6) 
      -- CP-element group 690: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1600_Update/$exit
      -- CP-element group 690: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1600_update_completed_
      -- CP-element group 690: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1602_Sample/req
      -- CP-element group 690: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1602_Sample/$entry
      -- CP-element group 690: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1602_sample_start_
      -- CP-element group 690: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1600_Update/ca
      -- 
    ca_3166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 690_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1600_inst_ack_1, ack => zeropad_CP_182_elements(690)); -- 
    req_3174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(690), ack => WPIPE_Zeropad_output_pipe_1602_inst_req_0); -- 
    -- CP-element group 691:  transition  input  output  bypass 
    -- CP-element group 691: predecessors 
    -- CP-element group 691: 	690 
    -- CP-element group 691: successors 
    -- CP-element group 691: 	692 
    -- CP-element group 691:  members (6) 
      -- CP-element group 691: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1602_Update/req
      -- CP-element group 691: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1602_Update/$entry
      -- CP-element group 691: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1602_Sample/ack
      -- CP-element group 691: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1602_Sample/$exit
      -- CP-element group 691: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1602_update_start_
      -- CP-element group 691: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1602_sample_completed_
      -- 
    ack_3175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 691_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1602_inst_ack_0, ack => zeropad_CP_182_elements(691)); -- 
    req_3179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(691), ack => WPIPE_Zeropad_output_pipe_1602_inst_req_1); -- 
    -- CP-element group 692:  transition  input  bypass 
    -- CP-element group 692: predecessors 
    -- CP-element group 692: 	691 
    -- CP-element group 692: successors 
    -- CP-element group 692: 	693 
    -- CP-element group 692:  members (3) 
      -- CP-element group 692: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1602_Update/ack
      -- CP-element group 692: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1602_Update/$exit
      -- CP-element group 692: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1602_update_completed_
      -- 
    ack_3180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 692_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1602_inst_ack_1, ack => zeropad_CP_182_elements(692)); -- 
    -- CP-element group 693:  join  transition  output  bypass 
    -- CP-element group 693: predecessors 
    -- CP-element group 693: 	688 
    -- CP-element group 693: 	692 
    -- CP-element group 693: successors 
    -- CP-element group 693: 	694 
    -- CP-element group 693:  members (3) 
      -- CP-element group 693: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1605_Sample/req
      -- CP-element group 693: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1605_Sample/$entry
      -- CP-element group 693: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1605_sample_start_
      -- 
    req_3188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(693), ack => WPIPE_Zeropad_output_pipe_1605_inst_req_0); -- 
    zeropad_cp_element_group_693: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_693"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(688) & zeropad_CP_182_elements(692);
      gj_zeropad_cp_element_group_693 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(693), clk => clk, reset => reset); --
    end block;
    -- CP-element group 694:  transition  input  output  bypass 
    -- CP-element group 694: predecessors 
    -- CP-element group 694: 	693 
    -- CP-element group 694: successors 
    -- CP-element group 694: 	695 
    -- CP-element group 694:  members (6) 
      -- CP-element group 694: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1605_Sample/$exit
      -- CP-element group 694: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1605_Sample/ack
      -- CP-element group 694: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1605_Update/$entry
      -- CP-element group 694: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1605_Update/req
      -- CP-element group 694: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1605_update_start_
      -- CP-element group 694: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1605_sample_completed_
      -- 
    ack_3189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 694_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1605_inst_ack_0, ack => zeropad_CP_182_elements(694)); -- 
    req_3193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(694), ack => WPIPE_Zeropad_output_pipe_1605_inst_req_1); -- 
    -- CP-element group 695:  transition  input  bypass 
    -- CP-element group 695: predecessors 
    -- CP-element group 695: 	694 
    -- CP-element group 695: successors 
    -- CP-element group 695: 	696 
    -- CP-element group 695:  members (3) 
      -- CP-element group 695: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1605_Update/$exit
      -- CP-element group 695: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1605_Update/ack
      -- CP-element group 695: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1605_update_completed_
      -- 
    ack_3194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 695_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1605_inst_ack_1, ack => zeropad_CP_182_elements(695)); -- 
    -- CP-element group 696:  join  transition  output  bypass 
    -- CP-element group 696: predecessors 
    -- CP-element group 696: 	686 
    -- CP-element group 696: 	695 
    -- CP-element group 696: successors 
    -- CP-element group 696: 	697 
    -- CP-element group 696:  members (3) 
      -- CP-element group 696: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1608_Sample/req
      -- CP-element group 696: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1608_sample_start_
      -- CP-element group 696: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1608_Sample/$entry
      -- 
    req_3202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(696), ack => WPIPE_Zeropad_output_pipe_1608_inst_req_0); -- 
    zeropad_cp_element_group_696: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_696"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(686) & zeropad_CP_182_elements(695);
      gj_zeropad_cp_element_group_696 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(696), clk => clk, reset => reset); --
    end block;
    -- CP-element group 697:  transition  input  output  bypass 
    -- CP-element group 697: predecessors 
    -- CP-element group 697: 	696 
    -- CP-element group 697: successors 
    -- CP-element group 697: 	698 
    -- CP-element group 697:  members (6) 
      -- CP-element group 697: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1608_Sample/$exit
      -- CP-element group 697: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1608_sample_completed_
      -- CP-element group 697: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1608_Update/req
      -- CP-element group 697: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1608_update_start_
      -- CP-element group 697: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1608_Update/$entry
      -- CP-element group 697: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1608_Sample/ack
      -- 
    ack_3203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 697_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1608_inst_ack_0, ack => zeropad_CP_182_elements(697)); -- 
    req_3207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(697), ack => WPIPE_Zeropad_output_pipe_1608_inst_req_1); -- 
    -- CP-element group 698:  transition  input  bypass 
    -- CP-element group 698: predecessors 
    -- CP-element group 698: 	697 
    -- CP-element group 698: successors 
    -- CP-element group 698: 	699 
    -- CP-element group 698:  members (3) 
      -- CP-element group 698: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1608_update_completed_
      -- CP-element group 698: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1608_Update/ack
      -- CP-element group 698: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1608_Update/$exit
      -- 
    ack_3208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 698_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1608_inst_ack_1, ack => zeropad_CP_182_elements(698)); -- 
    -- CP-element group 699:  join  transition  output  bypass 
    -- CP-element group 699: predecessors 
    -- CP-element group 699: 	684 
    -- CP-element group 699: 	698 
    -- CP-element group 699: successors 
    -- CP-element group 699: 	700 
    -- CP-element group 699:  members (3) 
      -- CP-element group 699: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1611_sample_start_
      -- CP-element group 699: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1611_Sample/req
      -- CP-element group 699: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1611_Sample/$entry
      -- 
    req_3216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(699), ack => WPIPE_Zeropad_output_pipe_1611_inst_req_0); -- 
    zeropad_cp_element_group_699: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_699"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(684) & zeropad_CP_182_elements(698);
      gj_zeropad_cp_element_group_699 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(699), clk => clk, reset => reset); --
    end block;
    -- CP-element group 700:  transition  input  output  bypass 
    -- CP-element group 700: predecessors 
    -- CP-element group 700: 	699 
    -- CP-element group 700: successors 
    -- CP-element group 700: 	701 
    -- CP-element group 700:  members (6) 
      -- CP-element group 700: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1611_update_start_
      -- CP-element group 700: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1611_sample_completed_
      -- CP-element group 700: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1611_Sample/ack
      -- CP-element group 700: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1611_Sample/$exit
      -- CP-element group 700: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1611_Update/$entry
      -- CP-element group 700: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1611_Update/req
      -- 
    ack_3217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 700_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1611_inst_ack_0, ack => zeropad_CP_182_elements(700)); -- 
    req_3221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(700), ack => WPIPE_Zeropad_output_pipe_1611_inst_req_1); -- 
    -- CP-element group 701:  transition  input  bypass 
    -- CP-element group 701: predecessors 
    -- CP-element group 701: 	700 
    -- CP-element group 701: successors 
    -- CP-element group 701: 	702 
    -- CP-element group 701:  members (3) 
      -- CP-element group 701: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1611_Update/ack
      -- CP-element group 701: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1611_update_completed_
      -- CP-element group 701: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1611_Update/$exit
      -- 
    ack_3222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 701_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1611_inst_ack_1, ack => zeropad_CP_182_elements(701)); -- 
    -- CP-element group 702:  join  transition  output  bypass 
    -- CP-element group 702: predecessors 
    -- CP-element group 702: 	682 
    -- CP-element group 702: 	701 
    -- CP-element group 702: successors 
    -- CP-element group 702: 	703 
    -- CP-element group 702:  members (3) 
      -- CP-element group 702: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1614_sample_start_
      -- CP-element group 702: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1614_Sample/$entry
      -- CP-element group 702: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1614_Sample/req
      -- 
    req_3230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(702), ack => WPIPE_Zeropad_output_pipe_1614_inst_req_0); -- 
    zeropad_cp_element_group_702: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_702"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(682) & zeropad_CP_182_elements(701);
      gj_zeropad_cp_element_group_702 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(702), clk => clk, reset => reset); --
    end block;
    -- CP-element group 703:  transition  input  output  bypass 
    -- CP-element group 703: predecessors 
    -- CP-element group 703: 	702 
    -- CP-element group 703: successors 
    -- CP-element group 703: 	704 
    -- CP-element group 703:  members (6) 
      -- CP-element group 703: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1614_Sample/ack
      -- CP-element group 703: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1614_Update/req
      -- CP-element group 703: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1614_Sample/$exit
      -- CP-element group 703: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1614_update_start_
      -- CP-element group 703: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1614_Update/$entry
      -- CP-element group 703: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1614_sample_completed_
      -- 
    ack_3231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 703_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1614_inst_ack_0, ack => zeropad_CP_182_elements(703)); -- 
    req_3235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(703), ack => WPIPE_Zeropad_output_pipe_1614_inst_req_1); -- 
    -- CP-element group 704:  transition  input  bypass 
    -- CP-element group 704: predecessors 
    -- CP-element group 704: 	703 
    -- CP-element group 704: successors 
    -- CP-element group 704: 	705 
    -- CP-element group 704:  members (3) 
      -- CP-element group 704: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1614_Update/ack
      -- CP-element group 704: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1614_update_completed_
      -- CP-element group 704: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1614_Update/$exit
      -- 
    ack_3236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 704_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1614_inst_ack_1, ack => zeropad_CP_182_elements(704)); -- 
    -- CP-element group 705:  join  transition  output  bypass 
    -- CP-element group 705: predecessors 
    -- CP-element group 705: 	680 
    -- CP-element group 705: 	704 
    -- CP-element group 705: successors 
    -- CP-element group 705: 	706 
    -- CP-element group 705:  members (3) 
      -- CP-element group 705: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1617_Sample/$entry
      -- CP-element group 705: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1617_Sample/req
      -- CP-element group 705: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1617_sample_start_
      -- 
    req_3244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(705), ack => WPIPE_Zeropad_output_pipe_1617_inst_req_0); -- 
    zeropad_cp_element_group_705: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_705"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(680) & zeropad_CP_182_elements(704);
      gj_zeropad_cp_element_group_705 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(705), clk => clk, reset => reset); --
    end block;
    -- CP-element group 706:  transition  input  output  bypass 
    -- CP-element group 706: predecessors 
    -- CP-element group 706: 	705 
    -- CP-element group 706: successors 
    -- CP-element group 706: 	707 
    -- CP-element group 706:  members (6) 
      -- CP-element group 706: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1617_update_start_
      -- CP-element group 706: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1617_sample_completed_
      -- CP-element group 706: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1617_Sample/ack
      -- CP-element group 706: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1617_Update/req
      -- CP-element group 706: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1617_Update/$entry
      -- CP-element group 706: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1617_Sample/$exit
      -- 
    ack_3245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 706_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1617_inst_ack_0, ack => zeropad_CP_182_elements(706)); -- 
    req_3249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(706), ack => WPIPE_Zeropad_output_pipe_1617_inst_req_1); -- 
    -- CP-element group 707:  transition  input  bypass 
    -- CP-element group 707: predecessors 
    -- CP-element group 707: 	706 
    -- CP-element group 707: successors 
    -- CP-element group 707: 	708 
    -- CP-element group 707:  members (3) 
      -- CP-element group 707: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1617_Update/ack
      -- CP-element group 707: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1617_Update/$exit
      -- CP-element group 707: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1617_update_completed_
      -- 
    ack_3250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 707_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1617_inst_ack_1, ack => zeropad_CP_182_elements(707)); -- 
    -- CP-element group 708:  join  transition  output  bypass 
    -- CP-element group 708: predecessors 
    -- CP-element group 708: 	678 
    -- CP-element group 708: 	707 
    -- CP-element group 708: successors 
    -- CP-element group 708: 	709 
    -- CP-element group 708:  members (3) 
      -- CP-element group 708: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1620_sample_start_
      -- CP-element group 708: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1620_Sample/$entry
      -- CP-element group 708: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1620_Sample/req
      -- 
    req_3258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(708), ack => WPIPE_Zeropad_output_pipe_1620_inst_req_0); -- 
    zeropad_cp_element_group_708: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_708"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(678) & zeropad_CP_182_elements(707);
      gj_zeropad_cp_element_group_708 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(708), clk => clk, reset => reset); --
    end block;
    -- CP-element group 709:  transition  input  output  bypass 
    -- CP-element group 709: predecessors 
    -- CP-element group 709: 	708 
    -- CP-element group 709: successors 
    -- CP-element group 709: 	710 
    -- CP-element group 709:  members (6) 
      -- CP-element group 709: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1620_sample_completed_
      -- CP-element group 709: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1620_update_start_
      -- CP-element group 709: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1620_Sample/$exit
      -- CP-element group 709: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1620_Sample/ack
      -- CP-element group 709: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1620_Update/$entry
      -- CP-element group 709: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1620_Update/req
      -- 
    ack_3259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 709_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1620_inst_ack_0, ack => zeropad_CP_182_elements(709)); -- 
    req_3263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(709), ack => WPIPE_Zeropad_output_pipe_1620_inst_req_1); -- 
    -- CP-element group 710:  transition  input  bypass 
    -- CP-element group 710: predecessors 
    -- CP-element group 710: 	709 
    -- CP-element group 710: successors 
    -- CP-element group 710: 	711 
    -- CP-element group 710:  members (3) 
      -- CP-element group 710: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1620_update_completed_
      -- CP-element group 710: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1620_Update/$exit
      -- CP-element group 710: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1620_Update/ack
      -- 
    ack_3264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 710_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1620_inst_ack_1, ack => zeropad_CP_182_elements(710)); -- 
    -- CP-element group 711:  join  transition  output  bypass 
    -- CP-element group 711: predecessors 
    -- CP-element group 711: 	676 
    -- CP-element group 711: 	710 
    -- CP-element group 711: successors 
    -- CP-element group 711: 	712 
    -- CP-element group 711:  members (3) 
      -- CP-element group 711: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1623_sample_start_
      -- CP-element group 711: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1623_Sample/$entry
      -- CP-element group 711: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1623_Sample/req
      -- 
    req_3272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(711), ack => WPIPE_Zeropad_output_pipe_1623_inst_req_0); -- 
    zeropad_cp_element_group_711: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_711"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(676) & zeropad_CP_182_elements(710);
      gj_zeropad_cp_element_group_711 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(711), clk => clk, reset => reset); --
    end block;
    -- CP-element group 712:  transition  input  output  bypass 
    -- CP-element group 712: predecessors 
    -- CP-element group 712: 	711 
    -- CP-element group 712: successors 
    -- CP-element group 712: 	713 
    -- CP-element group 712:  members (6) 
      -- CP-element group 712: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1623_sample_completed_
      -- CP-element group 712: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1623_update_start_
      -- CP-element group 712: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1623_Sample/$exit
      -- CP-element group 712: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1623_Sample/ack
      -- CP-element group 712: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1623_Update/$entry
      -- CP-element group 712: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1623_Update/req
      -- 
    ack_3273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 712_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1623_inst_ack_0, ack => zeropad_CP_182_elements(712)); -- 
    req_3277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(712), ack => WPIPE_Zeropad_output_pipe_1623_inst_req_1); -- 
    -- CP-element group 713:  transition  input  bypass 
    -- CP-element group 713: predecessors 
    -- CP-element group 713: 	712 
    -- CP-element group 713: successors 
    -- CP-element group 713: 	714 
    -- CP-element group 713:  members (3) 
      -- CP-element group 713: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1623_update_completed_
      -- CP-element group 713: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1623_Update/$exit
      -- CP-element group 713: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/WPIPE_Zeropad_output_pipe_1623_Update/ack
      -- 
    ack_3278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 713_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Zeropad_output_pipe_1623_inst_ack_1, ack => zeropad_CP_182_elements(713)); -- 
    -- CP-element group 714:  branch  join  transition  place  output  bypass 
    -- CP-element group 714: predecessors 
    -- CP-element group 714: 	669 
    -- CP-element group 714: 	713 
    -- CP-element group 714: successors 
    -- CP-element group 714: 	715 
    -- CP-element group 714: 	716 
    -- CP-element group 714:  members (10) 
      -- CP-element group 714: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636__exit__
      -- CP-element group 714: 	 branch_block_stmt_43/if_stmt_1637__entry__
      -- CP-element group 714: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/$exit
      -- CP-element group 714: 	 branch_block_stmt_43/if_stmt_1637_dead_link/$entry
      -- CP-element group 714: 	 branch_block_stmt_43/if_stmt_1637_eval_test/$entry
      -- CP-element group 714: 	 branch_block_stmt_43/if_stmt_1637_eval_test/$exit
      -- CP-element group 714: 	 branch_block_stmt_43/if_stmt_1637_eval_test/branch_req
      -- CP-element group 714: 	 branch_block_stmt_43/R_exitcond7_1638_place
      -- CP-element group 714: 	 branch_block_stmt_43/if_stmt_1637_if_link/$entry
      -- CP-element group 714: 	 branch_block_stmt_43/if_stmt_1637_else_link/$entry
      -- 
    branch_req_3286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(714), ack => if_stmt_1637_branch_req_0); -- 
    zeropad_cp_element_group_714: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_714"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(669) & zeropad_CP_182_elements(713);
      gj_zeropad_cp_element_group_714 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(714), clk => clk, reset => reset); --
    end block;
    -- CP-element group 715:  merge  transition  place  input  bypass 
    -- CP-element group 715: predecessors 
    -- CP-element group 715: 	714 
    -- CP-element group 715: successors 
    -- CP-element group 715: 	740 
    -- CP-element group 715:  members (13) 
      -- CP-element group 715: 	 branch_block_stmt_43/merge_stmt_1643__exit__
      -- CP-element group 715: 	 branch_block_stmt_43/forx_xend443x_xloopexit_forx_xend443
      -- CP-element group 715: 	 branch_block_stmt_43/if_stmt_1637_if_link/$exit
      -- CP-element group 715: 	 branch_block_stmt_43/if_stmt_1637_if_link/if_choice_transition
      -- CP-element group 715: 	 branch_block_stmt_43/forx_xbody371_forx_xend443x_xloopexit
      -- CP-element group 715: 	 branch_block_stmt_43/forx_xbody371_forx_xend443x_xloopexit_PhiReq/$entry
      -- CP-element group 715: 	 branch_block_stmt_43/forx_xbody371_forx_xend443x_xloopexit_PhiReq/$exit
      -- CP-element group 715: 	 branch_block_stmt_43/merge_stmt_1643_PhiReqMerge
      -- CP-element group 715: 	 branch_block_stmt_43/merge_stmt_1643_PhiAck/$entry
      -- CP-element group 715: 	 branch_block_stmt_43/merge_stmt_1643_PhiAck/$exit
      -- CP-element group 715: 	 branch_block_stmt_43/merge_stmt_1643_PhiAck/dummy
      -- CP-element group 715: 	 branch_block_stmt_43/forx_xend443x_xloopexit_forx_xend443_PhiReq/$entry
      -- CP-element group 715: 	 branch_block_stmt_43/forx_xend443x_xloopexit_forx_xend443_PhiReq/$exit
      -- 
    if_choice_transition_3291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 715_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1637_branch_ack_1, ack => zeropad_CP_182_elements(715)); -- 
    -- CP-element group 716:  fork  transition  place  input  output  bypass 
    -- CP-element group 716: predecessors 
    -- CP-element group 716: 	714 
    -- CP-element group 716: successors 
    -- CP-element group 716: 	735 
    -- CP-element group 716: 	736 
    -- CP-element group 716:  members (12) 
      -- CP-element group 716: 	 branch_block_stmt_43/if_stmt_1637_else_link/$exit
      -- CP-element group 716: 	 branch_block_stmt_43/if_stmt_1637_else_link/else_choice_transition
      -- CP-element group 716: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371
      -- CP-element group 716: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/$entry
      -- CP-element group 716: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1507/$entry
      -- CP-element group 716: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/$entry
      -- CP-element group 716: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1513/$entry
      -- CP-element group 716: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1513/SplitProtocol/$entry
      -- CP-element group 716: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1513/SplitProtocol/Sample/$entry
      -- CP-element group 716: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1513/SplitProtocol/Sample/rr
      -- CP-element group 716: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1513/SplitProtocol/Update/$entry
      -- CP-element group 716: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1513/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 716_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1637_branch_ack_0, ack => zeropad_CP_182_elements(716)); -- 
    rr_3483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(716), ack => type_cast_1513_inst_req_0); -- 
    cr_3488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(716), ack => type_cast_1513_inst_req_1); -- 
    -- CP-element group 717:  transition  output  delay-element  bypass 
    -- CP-element group 717: predecessors 
    -- CP-element group 717: 	57 
    -- CP-element group 717: successors 
    -- CP-element group 717: 	721 
    -- CP-element group 717:  members (5) 
      -- CP-element group 717: 	 branch_block_stmt_43/bbx_xnph464_forx_xbody_PhiReq/$exit
      -- CP-element group 717: 	 branch_block_stmt_43/bbx_xnph464_forx_xbody_PhiReq/phi_stmt_269/$exit
      -- CP-element group 717: 	 branch_block_stmt_43/bbx_xnph464_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_sources/$exit
      -- CP-element group 717: 	 branch_block_stmt_43/bbx_xnph464_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_273_konst_delay_trans
      -- CP-element group 717: 	 branch_block_stmt_43/bbx_xnph464_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_req
      -- 
    phi_stmt_269_req_3320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_269_req_3320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(717), ack => phi_stmt_269_req_0); -- 
    -- Element group zeropad_CP_182_elements(717) is a control-delay.
    cp_element_717_delay: control_delay_element  generic map(name => " 717_delay", delay_value => 1)  port map(req => zeropad_CP_182_elements(57), ack => zeropad_CP_182_elements(717), clk => clk, reset =>reset);
    -- CP-element group 718:  transition  input  bypass 
    -- CP-element group 718: predecessors 
    -- CP-element group 718: 	100 
    -- CP-element group 718: successors 
    -- CP-element group 718: 	720 
    -- CP-element group 718:  members (2) 
      -- CP-element group 718: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_275/SplitProtocol/Sample/$exit
      -- CP-element group 718: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_275/SplitProtocol/Sample/ra
      -- 
    ra_3340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 718_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_275_inst_ack_0, ack => zeropad_CP_182_elements(718)); -- 
    -- CP-element group 719:  transition  input  bypass 
    -- CP-element group 719: predecessors 
    -- CP-element group 719: 	100 
    -- CP-element group 719: successors 
    -- CP-element group 719: 	720 
    -- CP-element group 719:  members (2) 
      -- CP-element group 719: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_275/SplitProtocol/Update/$exit
      -- CP-element group 719: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_275/SplitProtocol/Update/ca
      -- 
    ca_3345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 719_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_275_inst_ack_1, ack => zeropad_CP_182_elements(719)); -- 
    -- CP-element group 720:  join  transition  output  bypass 
    -- CP-element group 720: predecessors 
    -- CP-element group 720: 	718 
    -- CP-element group 720: 	719 
    -- CP-element group 720: successors 
    -- CP-element group 720: 	721 
    -- CP-element group 720:  members (6) 
      -- CP-element group 720: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 720: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/phi_stmt_269/$exit
      -- CP-element group 720: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_sources/$exit
      -- CP-element group 720: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_275/$exit
      -- CP-element group 720: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_sources/type_cast_275/SplitProtocol/$exit
      -- CP-element group 720: 	 branch_block_stmt_43/forx_xbody_forx_xbody_PhiReq/phi_stmt_269/phi_stmt_269_req
      -- 
    phi_stmt_269_req_3346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_269_req_3346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(720), ack => phi_stmt_269_req_1); -- 
    zeropad_cp_element_group_720: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_720"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(718) & zeropad_CP_182_elements(719);
      gj_zeropad_cp_element_group_720 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(720), clk => clk, reset => reset); --
    end block;
    -- CP-element group 721:  merge  transition  place  bypass 
    -- CP-element group 721: predecessors 
    -- CP-element group 721: 	717 
    -- CP-element group 721: 	720 
    -- CP-element group 721: successors 
    -- CP-element group 721: 	722 
    -- CP-element group 721:  members (2) 
      -- CP-element group 721: 	 branch_block_stmt_43/merge_stmt_268_PhiReqMerge
      -- CP-element group 721: 	 branch_block_stmt_43/merge_stmt_268_PhiAck/$entry
      -- 
    zeropad_CP_182_elements(721) <= OrReduce(zeropad_CP_182_elements(717) & zeropad_CP_182_elements(720));
    -- CP-element group 722:  fork  transition  place  input  output  bypass 
    -- CP-element group 722: predecessors 
    -- CP-element group 722: 	721 
    -- CP-element group 722: successors 
    -- CP-element group 722: 	59 
    -- CP-element group 722: 	60 
    -- CP-element group 722: 	62 
    -- CP-element group 722: 	63 
    -- CP-element group 722: 	66 
    -- CP-element group 722: 	70 
    -- CP-element group 722: 	74 
    -- CP-element group 722: 	78 
    -- CP-element group 722: 	82 
    -- CP-element group 722: 	86 
    -- CP-element group 722: 	90 
    -- CP-element group 722: 	94 
    -- CP-element group 722: 	97 
    -- CP-element group 722:  members (56) 
      -- CP-element group 722: 	 branch_block_stmt_43/merge_stmt_268__exit__
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433__entry__
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/addr_of_284_complete/$entry
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/addr_of_284_complete/req
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_287_sample_start_
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_287_Sample/$entry
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/RPIPE_Zeropad_input_pipe_287_Sample/rr
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/$entry
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/addr_of_284_update_start_
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_index_resized_2
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_index_scaled_2
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_index_computed_2
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_index_resize_2/$entry
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_index_resize_2/$exit
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_index_resize_2/index_resize_req
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_index_resize_2/index_resize_ack
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_index_scale_2/$entry
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_index_scale_2/$exit
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_index_scale_2/scale_rename_req
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_index_scale_2/scale_rename_ack
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_final_index_sum_regn_update_start
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_final_index_sum_regn_Sample/$entry
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_final_index_sum_regn_Sample/req
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_final_index_sum_regn_Update/$entry
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/array_obj_ref_283_final_index_sum_regn_Update/req
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_291_update_start_
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_291_Update/$entry
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_291_Update/cr
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_304_update_start_
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_304_Update/$entry
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_304_Update/cr
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_322_update_start_
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_322_Update/$entry
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_322_Update/cr
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_340_update_start_
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_340_Update/$entry
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_340_Update/cr
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_358_update_start_
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_358_Update/$entry
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_358_Update/cr
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_376_update_start_
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_376_Update/$entry
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_376_Update/cr
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_394_update_start_
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_394_Update/$entry
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_394_Update/cr
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_412_update_start_
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_412_Update/$entry
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/type_cast_412_Update/cr
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_update_start_
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Update/$entry
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Update/word_access_complete/$entry
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Update/word_access_complete/word_0/$entry
      -- CP-element group 722: 	 branch_block_stmt_43/assign_stmt_285_to_assign_stmt_433/ptr_deref_420_Update/word_access_complete/word_0/cr
      -- CP-element group 722: 	 branch_block_stmt_43/merge_stmt_268_PhiAck/$exit
      -- CP-element group 722: 	 branch_block_stmt_43/merge_stmt_268_PhiAck/phi_stmt_269_ack
      -- 
    phi_stmt_269_ack_3351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 722_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_269_ack_0, ack => zeropad_CP_182_elements(722)); -- 
    req_680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(722), ack => addr_of_284_final_reg_req_1); -- 
    rr_689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(722), ack => RPIPE_Zeropad_input_pipe_287_inst_req_0); -- 
    req_660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(722), ack => array_obj_ref_283_index_offset_req_0); -- 
    req_665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(722), ack => array_obj_ref_283_index_offset_req_1); -- 
    cr_708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(722), ack => type_cast_291_inst_req_1); -- 
    cr_736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(722), ack => type_cast_304_inst_req_1); -- 
    cr_764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(722), ack => type_cast_322_inst_req_1); -- 
    cr_792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(722), ack => type_cast_340_inst_req_1); -- 
    cr_820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(722), ack => type_cast_358_inst_req_1); -- 
    cr_848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(722), ack => type_cast_376_inst_req_1); -- 
    cr_876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(722), ack => type_cast_394_inst_req_1); -- 
    cr_904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(722), ack => type_cast_412_inst_req_1); -- 
    cr_954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(722), ack => ptr_deref_420_store_0_req_1); -- 
    -- CP-element group 723:  merge  fork  transition  place  output  bypass 
    -- CP-element group 723: predecessors 
    -- CP-element group 723: 	58 
    -- CP-element group 723: 	99 
    -- CP-element group 723: successors 
    -- CP-element group 723: 	101 
    -- CP-element group 723: 	102 
    -- CP-element group 723:  members (13) 
      -- CP-element group 723: 	 branch_block_stmt_43/merge_stmt_442__exit__
      -- CP-element group 723: 	 branch_block_stmt_43/call_stmt_445__entry__
      -- CP-element group 723: 	 branch_block_stmt_43/call_stmt_445/$entry
      -- CP-element group 723: 	 branch_block_stmt_43/call_stmt_445/call_stmt_445_sample_start_
      -- CP-element group 723: 	 branch_block_stmt_43/call_stmt_445/call_stmt_445_update_start_
      -- CP-element group 723: 	 branch_block_stmt_43/call_stmt_445/call_stmt_445_Sample/$entry
      -- CP-element group 723: 	 branch_block_stmt_43/call_stmt_445/call_stmt_445_Sample/crr
      -- CP-element group 723: 	 branch_block_stmt_43/call_stmt_445/call_stmt_445_Update/$entry
      -- CP-element group 723: 	 branch_block_stmt_43/call_stmt_445/call_stmt_445_Update/ccr
      -- CP-element group 723: 	 branch_block_stmt_43/merge_stmt_442_PhiReqMerge
      -- CP-element group 723: 	 branch_block_stmt_43/merge_stmt_442_PhiAck/$entry
      -- CP-element group 723: 	 branch_block_stmt_43/merge_stmt_442_PhiAck/$exit
      -- CP-element group 723: 	 branch_block_stmt_43/merge_stmt_442_PhiAck/dummy
      -- 
    crr_985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(723), ack => call_stmt_445_call_req_0); -- 
    ccr_990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(723), ack => call_stmt_445_call_req_1); -- 
    zeropad_CP_182_elements(723) <= OrReduce(zeropad_CP_182_elements(58) & zeropad_CP_182_elements(99));
    -- CP-element group 724:  transition  input  bypass 
    -- CP-element group 724: predecessors 
    -- CP-element group 724: 	104 
    -- CP-element group 724: successors 
    -- CP-element group 724: 	726 
    -- CP-element group 724:  members (2) 
      -- CP-element group 724: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_539/phi_stmt_539_sources/type_cast_542/SplitProtocol/Sample/$exit
      -- CP-element group 724: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_539/phi_stmt_539_sources/type_cast_542/SplitProtocol/Sample/ra
      -- 
    ra_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 724_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_542_inst_ack_0, ack => zeropad_CP_182_elements(724)); -- 
    -- CP-element group 725:  transition  input  bypass 
    -- CP-element group 725: predecessors 
    -- CP-element group 725: 	104 
    -- CP-element group 725: successors 
    -- CP-element group 725: 	726 
    -- CP-element group 725:  members (2) 
      -- CP-element group 725: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_539/phi_stmt_539_sources/type_cast_542/SplitProtocol/Update/$exit
      -- CP-element group 725: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_539/phi_stmt_539_sources/type_cast_542/SplitProtocol/Update/ca
      -- 
    ca_3399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 725_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_542_inst_ack_1, ack => zeropad_CP_182_elements(725)); -- 
    -- CP-element group 726:  join  transition  output  bypass 
    -- CP-element group 726: predecessors 
    -- CP-element group 726: 	724 
    -- CP-element group 726: 	725 
    -- CP-element group 726: successors 
    -- CP-element group 726: 	730 
    -- CP-element group 726:  members (5) 
      -- CP-element group 726: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_539/$exit
      -- CP-element group 726: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_539/phi_stmt_539_sources/$exit
      -- CP-element group 726: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_539/phi_stmt_539_sources/type_cast_542/$exit
      -- CP-element group 726: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_539/phi_stmt_539_sources/type_cast_542/SplitProtocol/$exit
      -- CP-element group 726: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_539/phi_stmt_539_req
      -- 
    phi_stmt_539_req_3400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_539_req_3400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(726), ack => phi_stmt_539_req_0); -- 
    zeropad_cp_element_group_726: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_726"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(724) & zeropad_CP_182_elements(725);
      gj_zeropad_cp_element_group_726 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(726), clk => clk, reset => reset); --
    end block;
    -- CP-element group 727:  transition  input  bypass 
    -- CP-element group 727: predecessors 
    -- CP-element group 727: 	104 
    -- CP-element group 727: successors 
    -- CP-element group 727: 	729 
    -- CP-element group 727:  members (2) 
      -- CP-element group 727: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_586/SplitProtocol/Sample/$exit
      -- CP-element group 727: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_586/SplitProtocol/Sample/ra
      -- 
    ra_3417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 727_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_586_inst_ack_0, ack => zeropad_CP_182_elements(727)); -- 
    -- CP-element group 728:  transition  input  bypass 
    -- CP-element group 728: predecessors 
    -- CP-element group 728: 	104 
    -- CP-element group 728: successors 
    -- CP-element group 728: 	729 
    -- CP-element group 728:  members (2) 
      -- CP-element group 728: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_586/SplitProtocol/Update/$exit
      -- CP-element group 728: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_586/SplitProtocol/Update/ca
      -- 
    ca_3422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 728_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_586_inst_ack_1, ack => zeropad_CP_182_elements(728)); -- 
    -- CP-element group 729:  join  transition  output  bypass 
    -- CP-element group 729: predecessors 
    -- CP-element group 729: 	727 
    -- CP-element group 729: 	728 
    -- CP-element group 729: successors 
    -- CP-element group 729: 	730 
    -- CP-element group 729:  members (5) 
      -- CP-element group 729: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_583/$exit
      -- CP-element group 729: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_583/phi_stmt_583_sources/$exit
      -- CP-element group 729: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_586/$exit
      -- CP-element group 729: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_583/phi_stmt_583_sources/type_cast_586/SplitProtocol/$exit
      -- CP-element group 729: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/phi_stmt_583/phi_stmt_583_req
      -- 
    phi_stmt_583_req_3423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_583_req_3423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(729), ack => phi_stmt_583_req_0); -- 
    zeropad_cp_element_group_729: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_729"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(727) & zeropad_CP_182_elements(728);
      gj_zeropad_cp_element_group_729 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(729), clk => clk, reset => reset); --
    end block;
    -- CP-element group 730:  join  fork  transition  place  bypass 
    -- CP-element group 730: predecessors 
    -- CP-element group 730: 	726 
    -- CP-element group 730: 	729 
    -- CP-element group 730: successors 
    -- CP-element group 730: 	731 
    -- CP-element group 730: 	732 
    -- CP-element group 730:  members (3) 
      -- CP-element group 730: 	 branch_block_stmt_43/forx_xend_whilex_xbody_PhiReq/$exit
      -- CP-element group 730: 	 branch_block_stmt_43/merge_stmt_533_PhiReqMerge
      -- CP-element group 730: 	 branch_block_stmt_43/merge_stmt_533_PhiAck/$entry
      -- 
    zeropad_cp_element_group_730: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_730"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(726) & zeropad_CP_182_elements(729);
      gj_zeropad_cp_element_group_730 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(730), clk => clk, reset => reset); --
    end block;
    -- CP-element group 731:  transition  input  bypass 
    -- CP-element group 731: predecessors 
    -- CP-element group 731: 	730 
    -- CP-element group 731: successors 
    -- CP-element group 731: 	733 
    -- CP-element group 731:  members (1) 
      -- CP-element group 731: 	 branch_block_stmt_43/merge_stmt_533_PhiAck/phi_stmt_539_ack
      -- 
    phi_stmt_539_ack_3428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 731_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_539_ack_0, ack => zeropad_CP_182_elements(731)); -- 
    -- CP-element group 732:  transition  input  bypass 
    -- CP-element group 732: predecessors 
    -- CP-element group 732: 	730 
    -- CP-element group 732: successors 
    -- CP-element group 732: 	733 
    -- CP-element group 732:  members (1) 
      -- CP-element group 732: 	 branch_block_stmt_43/merge_stmt_533_PhiAck/phi_stmt_583_ack
      -- 
    phi_stmt_583_ack_3429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 732_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_583_ack_0, ack => zeropad_CP_182_elements(732)); -- 
    -- CP-element group 733:  join  transition  place  bypass 
    -- CP-element group 733: predecessors 
    -- CP-element group 733: 	731 
    -- CP-element group 733: 	732 
    -- CP-element group 733: successors 
    -- CP-element group 733: 	105 
    -- CP-element group 733:  members (3) 
      -- CP-element group 733: 	 branch_block_stmt_43/merge_stmt_533__exit__
      -- CP-element group 733: 	 branch_block_stmt_43/do_while_stmt_588__entry__
      -- CP-element group 733: 	 branch_block_stmt_43/merge_stmt_533_PhiAck/$exit
      -- 
    zeropad_cp_element_group_733: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_733"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(731) & zeropad_CP_182_elements(732);
      gj_zeropad_cp_element_group_733 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(733), clk => clk, reset => reset); --
    end block;
    -- CP-element group 734:  transition  output  delay-element  bypass 
    -- CP-element group 734: predecessors 
    -- CP-element group 734: 	668 
    -- CP-element group 734: successors 
    -- CP-element group 734: 	738 
    -- CP-element group 734:  members (5) 
      -- CP-element group 734: 	 branch_block_stmt_43/bbx_xnph_forx_xbody371_PhiReq/$exit
      -- CP-element group 734: 	 branch_block_stmt_43/bbx_xnph_forx_xbody371_PhiReq/phi_stmt_1507/$exit
      -- CP-element group 734: 	 branch_block_stmt_43/bbx_xnph_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/$exit
      -- CP-element group 734: 	 branch_block_stmt_43/bbx_xnph_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1511_konst_delay_trans
      -- CP-element group 734: 	 branch_block_stmt_43/bbx_xnph_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_req
      -- 
    phi_stmt_1507_req_3464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1507_req_3464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(734), ack => phi_stmt_1507_req_0); -- 
    -- Element group zeropad_CP_182_elements(734) is a control-delay.
    cp_element_734_delay: control_delay_element  generic map(name => " 734_delay", delay_value => 1)  port map(req => zeropad_CP_182_elements(668), ack => zeropad_CP_182_elements(734), clk => clk, reset =>reset);
    -- CP-element group 735:  transition  input  bypass 
    -- CP-element group 735: predecessors 
    -- CP-element group 735: 	716 
    -- CP-element group 735: successors 
    -- CP-element group 735: 	737 
    -- CP-element group 735:  members (2) 
      -- CP-element group 735: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1513/SplitProtocol/Sample/$exit
      -- CP-element group 735: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1513/SplitProtocol/Sample/ra
      -- 
    ra_3484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 735_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1513_inst_ack_0, ack => zeropad_CP_182_elements(735)); -- 
    -- CP-element group 736:  transition  input  bypass 
    -- CP-element group 736: predecessors 
    -- CP-element group 736: 	716 
    -- CP-element group 736: successors 
    -- CP-element group 736: 	737 
    -- CP-element group 736:  members (2) 
      -- CP-element group 736: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1513/SplitProtocol/Update/$exit
      -- CP-element group 736: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1513/SplitProtocol/Update/ca
      -- 
    ca_3489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 736_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1513_inst_ack_1, ack => zeropad_CP_182_elements(736)); -- 
    -- CP-element group 737:  join  transition  output  bypass 
    -- CP-element group 737: predecessors 
    -- CP-element group 737: 	735 
    -- CP-element group 737: 	736 
    -- CP-element group 737: successors 
    -- CP-element group 737: 	738 
    -- CP-element group 737:  members (6) 
      -- CP-element group 737: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/$exit
      -- CP-element group 737: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1507/$exit
      -- CP-element group 737: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/$exit
      -- CP-element group 737: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1513/$exit
      -- CP-element group 737: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1513/SplitProtocol/$exit
      -- CP-element group 737: 	 branch_block_stmt_43/forx_xbody371_forx_xbody371_PhiReq/phi_stmt_1507/phi_stmt_1507_req
      -- 
    phi_stmt_1507_req_3490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1507_req_3490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(737), ack => phi_stmt_1507_req_1); -- 
    zeropad_cp_element_group_737: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "zeropad_cp_element_group_737"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad_CP_182_elements(735) & zeropad_CP_182_elements(736);
      gj_zeropad_cp_element_group_737 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad_CP_182_elements(737), clk => clk, reset => reset); --
    end block;
    -- CP-element group 738:  merge  transition  place  bypass 
    -- CP-element group 738: predecessors 
    -- CP-element group 738: 	734 
    -- CP-element group 738: 	737 
    -- CP-element group 738: successors 
    -- CP-element group 738: 	739 
    -- CP-element group 738:  members (2) 
      -- CP-element group 738: 	 branch_block_stmt_43/merge_stmt_1506_PhiReqMerge
      -- CP-element group 738: 	 branch_block_stmt_43/merge_stmt_1506_PhiAck/$entry
      -- 
    zeropad_CP_182_elements(738) <= OrReduce(zeropad_CP_182_elements(734) & zeropad_CP_182_elements(737));
    -- CP-element group 739:  fork  transition  place  input  output  bypass 
    -- CP-element group 739: predecessors 
    -- CP-element group 739: 	738 
    -- CP-element group 739: successors 
    -- CP-element group 739: 	669 
    -- CP-element group 739: 	670 
    -- CP-element group 739: 	672 
    -- CP-element group 739: 	674 
    -- CP-element group 739: 	676 
    -- CP-element group 739: 	678 
    -- CP-element group 739: 	680 
    -- CP-element group 739: 	682 
    -- CP-element group 739: 	684 
    -- CP-element group 739: 	686 
    -- CP-element group 739: 	688 
    -- CP-element group 739: 	690 
    -- CP-element group 739:  members (53) 
      -- CP-element group 739: 	 branch_block_stmt_43/merge_stmt_1506__exit__
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636__entry__
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1530_Update/$entry
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1530_Update/cr
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Update/$entry
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1590_update_start_
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1550_update_start_
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Update/word_access_complete/word_0/$entry
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_final_index_sum_regn_Sample/$entry
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_final_index_sum_regn_Update/$entry
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Update/word_access_complete/$entry
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1580_Update/cr
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_final_index_sum_regn_Sample/req
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_index_scale_2/scale_rename_ack
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1590_Update/$entry
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_final_index_sum_regn_update_start
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1540_Update/cr
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_Update/word_access_complete/word_0/cr
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1590_Update/cr
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_final_index_sum_regn_Update/req
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1550_Update/$entry
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1600_update_start_
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1550_Update/cr
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1540_update_start_
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/addr_of_1522_complete/$entry
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/addr_of_1522_complete/req
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1530_update_start_
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1600_Update/$entry
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1560_update_start_
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/ptr_deref_1526_update_start_
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_index_scale_2/scale_rename_req
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_index_scale_2/$exit
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1580_Update/$entry
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_index_scale_2/$entry
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_index_resize_2/index_resize_ack
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_index_resize_2/index_resize_req
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_index_resize_2/$exit
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_index_resize_2/$entry
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1580_update_start_
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_index_computed_2
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_index_scaled_2
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/array_obj_ref_1521_index_resized_2
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1540_Update/$entry
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1570_Update/cr
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1570_Update/$entry
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/addr_of_1522_update_start_
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1570_update_start_
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1600_Update/cr
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/$entry
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1560_Update/cr
      -- CP-element group 739: 	 branch_block_stmt_43/assign_stmt_1523_to_assign_stmt_1636/type_cast_1560_Update/$entry
      -- CP-element group 739: 	 branch_block_stmt_43/merge_stmt_1506_PhiAck/$exit
      -- CP-element group 739: 	 branch_block_stmt_43/merge_stmt_1506_PhiAck/phi_stmt_1507_ack
      -- 
    phi_stmt_1507_ack_3495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 739_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1507_ack_0, ack => zeropad_CP_182_elements(739)); -- 
    cr_3067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(739), ack => type_cast_1530_inst_req_1); -- 
    cr_3137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(739), ack => type_cast_1580_inst_req_1); -- 
    req_2983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(739), ack => array_obj_ref_1521_index_offset_req_0); -- 
    cr_3081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(739), ack => type_cast_1540_inst_req_1); -- 
    cr_3048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(739), ack => ptr_deref_1526_load_0_req_1); -- 
    cr_3151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(739), ack => type_cast_1590_inst_req_1); -- 
    req_2988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(739), ack => array_obj_ref_1521_index_offset_req_1); -- 
    cr_3095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(739), ack => type_cast_1550_inst_req_1); -- 
    req_3003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(739), ack => addr_of_1522_final_reg_req_1); -- 
    cr_3123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(739), ack => type_cast_1570_inst_req_1); -- 
    cr_3165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(739), ack => type_cast_1600_inst_req_1); -- 
    cr_3109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad_CP_182_elements(739), ack => type_cast_1560_inst_req_1); -- 
    -- CP-element group 740:  merge  transition  place  bypass 
    -- CP-element group 740: predecessors 
    -- CP-element group 740: 	663 
    -- CP-element group 740: 	715 
    -- CP-element group 740: successors 
    -- CP-element group 740:  members (16) 
      -- CP-element group 740: 	 $exit
      -- CP-element group 740: 	 branch_block_stmt_43/$exit
      -- CP-element group 740: 	 branch_block_stmt_43/branch_block_stmt_43__exit__
      -- CP-element group 740: 	 branch_block_stmt_43/merge_stmt_1645__exit__
      -- CP-element group 740: 	 branch_block_stmt_43/return__
      -- CP-element group 740: 	 branch_block_stmt_43/merge_stmt_1647__exit__
      -- CP-element group 740: 	 branch_block_stmt_43/merge_stmt_1645_PhiReqMerge
      -- CP-element group 740: 	 branch_block_stmt_43/merge_stmt_1645_PhiAck/$entry
      -- CP-element group 740: 	 branch_block_stmt_43/merge_stmt_1645_PhiAck/$exit
      -- CP-element group 740: 	 branch_block_stmt_43/merge_stmt_1645_PhiAck/dummy
      -- CP-element group 740: 	 branch_block_stmt_43/return___PhiReq/$entry
      -- CP-element group 740: 	 branch_block_stmt_43/return___PhiReq/$exit
      -- CP-element group 740: 	 branch_block_stmt_43/merge_stmt_1647_PhiReqMerge
      -- CP-element group 740: 	 branch_block_stmt_43/merge_stmt_1647_PhiAck/$entry
      -- CP-element group 740: 	 branch_block_stmt_43/merge_stmt_1647_PhiAck/$exit
      -- CP-element group 740: 	 branch_block_stmt_43/merge_stmt_1647_PhiAck/dummy
      -- 
    zeropad_CP_182_elements(740) <= OrReduce(zeropad_CP_182_elements(663) & zeropad_CP_182_elements(715));
    zeropad_do_while_stmt_588_terminator_2612: loop_terminator -- 
      generic map (name => " zeropad_do_while_stmt_588_terminator_2612", max_iterations_in_flight =>15) 
      port map(loop_body_exit => zeropad_CP_182_elements(109),loop_continue => zeropad_CP_182_elements(613),loop_terminate => zeropad_CP_182_elements(612),loop_back => zeropad_CP_182_elements(107),loop_exit => zeropad_CP_182_elements(106),clk => clk, reset => reset); -- 
    phi_stmt_590_phi_seq_1108_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_CP_182_elements(122);
      zeropad_CP_182_elements(127)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_CP_182_elements(131);
      zeropad_CP_182_elements(128)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_CP_182_elements(132);
      zeropad_CP_182_elements(123) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_CP_182_elements(124);
      zeropad_CP_182_elements(133)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_CP_182_elements(133);
      zeropad_CP_182_elements(134)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_CP_182_elements(135);
      zeropad_CP_182_elements(125) <= phi_mux_reqs(1);
      phi_stmt_590_phi_seq_1108 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_590_phi_seq_1108") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_CP_182_elements(114), 
          phi_sample_ack => zeropad_CP_182_elements(120), 
          phi_update_req => zeropad_CP_182_elements(116), 
          phi_update_ack => zeropad_CP_182_elements(121), 
          phi_mux_ack => zeropad_CP_182_elements(126), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_595_phi_seq_1162_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_CP_182_elements(143);
      zeropad_CP_182_elements(148)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_CP_182_elements(152);
      zeropad_CP_182_elements(149)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_CP_182_elements(153);
      zeropad_CP_182_elements(144) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_CP_182_elements(145);
      zeropad_CP_182_elements(154)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_CP_182_elements(156);
      zeropad_CP_182_elements(155)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_CP_182_elements(157);
      zeropad_CP_182_elements(146) <= phi_mux_reqs(1);
      phi_stmt_595_phi_seq_1162 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_595_phi_seq_1162") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_CP_182_elements(139), 
          phi_sample_ack => zeropad_CP_182_elements(140), 
          phi_update_req => zeropad_CP_182_elements(141), 
          phi_update_ack => zeropad_CP_182_elements(142), 
          phi_mux_ack => zeropad_CP_182_elements(147), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_600_phi_seq_1206_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_CP_182_elements(164);
      zeropad_CP_182_elements(169)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_CP_182_elements(173);
      zeropad_CP_182_elements(170)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_CP_182_elements(174);
      zeropad_CP_182_elements(165) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_CP_182_elements(166);
      zeropad_CP_182_elements(175)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_CP_182_elements(175);
      zeropad_CP_182_elements(176)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_CP_182_elements(177);
      zeropad_CP_182_elements(167) <= phi_mux_reqs(1);
      phi_stmt_600_phi_seq_1206 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_600_phi_seq_1206") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_CP_182_elements(160), 
          phi_sample_ack => zeropad_CP_182_elements(161), 
          phi_update_req => zeropad_CP_182_elements(162), 
          phi_update_ack => zeropad_CP_182_elements(163), 
          phi_mux_ack => zeropad_CP_182_elements(168), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_605_phi_seq_1250_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_CP_182_elements(185);
      zeropad_CP_182_elements(190)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_CP_182_elements(194);
      zeropad_CP_182_elements(191)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_CP_182_elements(195);
      zeropad_CP_182_elements(186) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_CP_182_elements(187);
      zeropad_CP_182_elements(196)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_CP_182_elements(196);
      zeropad_CP_182_elements(197)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_CP_182_elements(198);
      zeropad_CP_182_elements(188) <= phi_mux_reqs(1);
      phi_stmt_605_phi_seq_1250 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_605_phi_seq_1250") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_CP_182_elements(181), 
          phi_sample_ack => zeropad_CP_182_elements(182), 
          phi_update_req => zeropad_CP_182_elements(183), 
          phi_update_ack => zeropad_CP_182_elements(184), 
          phi_mux_ack => zeropad_CP_182_elements(189), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_610_phi_seq_1294_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_CP_182_elements(206);
      zeropad_CP_182_elements(211)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_CP_182_elements(215);
      zeropad_CP_182_elements(212)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_CP_182_elements(216);
      zeropad_CP_182_elements(207) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_CP_182_elements(208);
      zeropad_CP_182_elements(217)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_CP_182_elements(217);
      zeropad_CP_182_elements(218)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_CP_182_elements(219);
      zeropad_CP_182_elements(209) <= phi_mux_reqs(1);
      phi_stmt_610_phi_seq_1294 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_610_phi_seq_1294") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_CP_182_elements(202), 
          phi_sample_ack => zeropad_CP_182_elements(203), 
          phi_update_req => zeropad_CP_182_elements(204), 
          phi_update_ack => zeropad_CP_182_elements(205), 
          phi_mux_ack => zeropad_CP_182_elements(210), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_615_phi_seq_1338_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_CP_182_elements(227);
      zeropad_CP_182_elements(232)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_CP_182_elements(236);
      zeropad_CP_182_elements(233)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_CP_182_elements(237);
      zeropad_CP_182_elements(228) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_CP_182_elements(229);
      zeropad_CP_182_elements(238)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_CP_182_elements(238);
      zeropad_CP_182_elements(239)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_CP_182_elements(240);
      zeropad_CP_182_elements(230) <= phi_mux_reqs(1);
      phi_stmt_615_phi_seq_1338 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_615_phi_seq_1338") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_CP_182_elements(223), 
          phi_sample_ack => zeropad_CP_182_elements(224), 
          phi_update_req => zeropad_CP_182_elements(225), 
          phi_update_ack => zeropad_CP_182_elements(226), 
          phi_mux_ack => zeropad_CP_182_elements(231), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_620_phi_seq_1382_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_CP_182_elements(248);
      zeropad_CP_182_elements(253)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_CP_182_elements(257);
      zeropad_CP_182_elements(254)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_CP_182_elements(258);
      zeropad_CP_182_elements(249) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_CP_182_elements(250);
      zeropad_CP_182_elements(259)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_CP_182_elements(259);
      zeropad_CP_182_elements(260)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_CP_182_elements(261);
      zeropad_CP_182_elements(251) <= phi_mux_reqs(1);
      phi_stmt_620_phi_seq_1382 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_620_phi_seq_1382") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_CP_182_elements(244), 
          phi_sample_ack => zeropad_CP_182_elements(245), 
          phi_update_req => zeropad_CP_182_elements(246), 
          phi_update_ack => zeropad_CP_182_elements(247), 
          phi_mux_ack => zeropad_CP_182_elements(252), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_625_phi_seq_1426_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_CP_182_elements(269);
      zeropad_CP_182_elements(274)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_CP_182_elements(278);
      zeropad_CP_182_elements(275)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_CP_182_elements(279);
      zeropad_CP_182_elements(270) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_CP_182_elements(271);
      zeropad_CP_182_elements(280)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_CP_182_elements(280);
      zeropad_CP_182_elements(281)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_CP_182_elements(282);
      zeropad_CP_182_elements(272) <= phi_mux_reqs(1);
      phi_stmt_625_phi_seq_1426 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_625_phi_seq_1426") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_CP_182_elements(265), 
          phi_sample_ack => zeropad_CP_182_elements(266), 
          phi_update_req => zeropad_CP_182_elements(267), 
          phi_update_ack => zeropad_CP_182_elements(268), 
          phi_mux_ack => zeropad_CP_182_elements(273), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_630_phi_seq_1470_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_CP_182_elements(290);
      zeropad_CP_182_elements(295)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_CP_182_elements(299);
      zeropad_CP_182_elements(296)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_CP_182_elements(300);
      zeropad_CP_182_elements(291) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_CP_182_elements(292);
      zeropad_CP_182_elements(301)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_CP_182_elements(301);
      zeropad_CP_182_elements(302)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_CP_182_elements(303);
      zeropad_CP_182_elements(293) <= phi_mux_reqs(1);
      phi_stmt_630_phi_seq_1470 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_630_phi_seq_1470") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_CP_182_elements(286), 
          phi_sample_ack => zeropad_CP_182_elements(287), 
          phi_update_req => zeropad_CP_182_elements(288), 
          phi_update_ack => zeropad_CP_182_elements(289), 
          phi_mux_ack => zeropad_CP_182_elements(294), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_635_phi_seq_1514_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_CP_182_elements(311);
      zeropad_CP_182_elements(316)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_CP_182_elements(320);
      zeropad_CP_182_elements(317)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_CP_182_elements(321);
      zeropad_CP_182_elements(312) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_CP_182_elements(313);
      zeropad_CP_182_elements(322)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_CP_182_elements(322);
      zeropad_CP_182_elements(323)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_CP_182_elements(324);
      zeropad_CP_182_elements(314) <= phi_mux_reqs(1);
      phi_stmt_635_phi_seq_1514 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_635_phi_seq_1514") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_CP_182_elements(307), 
          phi_sample_ack => zeropad_CP_182_elements(308), 
          phi_update_req => zeropad_CP_182_elements(309), 
          phi_update_ack => zeropad_CP_182_elements(310), 
          phi_mux_ack => zeropad_CP_182_elements(315), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_640_phi_seq_1568_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad_CP_182_elements(332);
      zeropad_CP_182_elements(337)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad_CP_182_elements(341);
      zeropad_CP_182_elements(338)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad_CP_182_elements(342);
      zeropad_CP_182_elements(333) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad_CP_182_elements(334);
      zeropad_CP_182_elements(343)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad_CP_182_elements(345);
      zeropad_CP_182_elements(344)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad_CP_182_elements(346);
      zeropad_CP_182_elements(335) <= phi_mux_reqs(1);
      phi_stmt_640_phi_seq_1568 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_640_phi_seq_1568") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad_CP_182_elements(328), 
          phi_sample_ack => zeropad_CP_182_elements(329), 
          phi_update_req => zeropad_CP_182_elements(330), 
          phi_update_ack => zeropad_CP_182_elements(331), 
          phi_mux_ack => zeropad_CP_182_elements(336), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1060_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= zeropad_CP_182_elements(110);
        preds(1)  <= zeropad_CP_182_elements(111);
        entry_tmerge_1060 : transition_merge -- 
          generic map(name => " entry_tmerge_1060")
          port map (preds => preds, symbol_out => zeropad_CP_182_elements(112));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal MUX_1005_1005_delayed_3_0_1132 : std_logic_vector(31 downto 0);
    signal MUX_1028_wire : std_logic_vector(31 downto 0);
    signal MUX_1029_wire : std_logic_vector(31 downto 0);
    signal MUX_1220_wire : std_logic_vector(31 downto 0);
    signal MUX_1233_wire : std_logic_vector(7 downto 0);
    signal MUX_1246_wire : std_logic_vector(63 downto 0);
    signal MUX_815_815_delayed_12_0_843 : std_logic_vector(63 downto 0);
    signal MUX_817_wire : std_logic_vector(31 downto 0);
    signal MUX_830_wire : std_logic_vector(7 downto 0);
    signal MUX_957_957_delayed_12_0_1063 : std_logic_vector(63 downto 0);
    signal MUX_969_969_delayed_2_0_1082 : std_logic_vector(7 downto 0);
    signal MUX_981_981_delayed_2_0_1100 : std_logic_vector(31 downto 0);
    signal MUX_993_993_delayed_2_0_1114 : std_logic_vector(63 downto 0);
    signal NOT_u1_u1_1175_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1331_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_770_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_903_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_940_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_998_wire : std_logic_vector(0 downto 0);
    signal R_add182_788_resized : std_logic_vector(14 downto 0);
    signal R_add182_788_scaled : std_logic_vector(14 downto 0);
    signal R_add_outx_x1_1186_resized : std_logic_vector(14 downto 0);
    signal R_add_outx_x1_1186_scaled : std_logic_vector(14 downto 0);
    signal R_ix_x0463_282_resized : std_logic_vector(14 downto 0);
    signal R_ix_x0463_282_scaled : std_logic_vector(14 downto 0);
    signal R_ix_x1460_1520_resized : std_logic_vector(14 downto 0);
    signal R_ix_x1460_1520_scaled : std_logic_vector(14 downto 0);
    signal add103_382 : std_logic_vector(63 downto 0);
    signal add109_400 : std_logic_vector(63 downto 0);
    signal add115_418 : std_logic_vector(63 downto 0);
    signal add12_94 : std_logic_vector(31 downto 0);
    signal add144_473 : std_logic_vector(31 downto 0);
    signal add173_754 : std_logic_vector(63 downto 0);
    signal add182_782 : std_logic_vector(31 downto 0);
    signal add21_119 : std_logic_vector(31 downto 0);
    signal add234_903_delayed_1_0_977 : std_logic_vector(31 downto 0);
    signal add234_962 : std_logic_vector(31 downto 0);
    signal add234x_xtarget_out_offsetx_x1_987 : std_logic_vector(31 downto 0);
    signal add30_145 : std_logic_vector(15 downto 0);
    signal add39_170 : std_logic_vector(15 downto 0);
    signal add48_195 : std_logic_vector(31 downto 0);
    signal add79_310 : std_logic_vector(63 downto 0);
    signal add85_328 : std_logic_vector(63 downto 0);
    signal add91_346 : std_logic_vector(63 downto 0);
    signal add97_364 : std_logic_vector(63 downto 0);
    signal add_69 : std_logic_vector(31 downto 0);
    signal add_outx_x0_1222 : std_logic_vector(31 downto 0);
    signal add_outx_x1_1059_delayed_2_0_1197 : std_logic_vector(31 downto 0);
    signal add_outx_x1_605 : std_logic_vector(31 downto 0);
    signal add_outx_x1_at_entry_548 : std_logic_vector(31 downto 0);
    signal add_srcx_x0452_1106 : std_logic_vector(31 downto 0);
    signal add_srcx_x0x_xph_819 : std_logic_vector(31 downto 0);
    signal add_srcx_x1_590 : std_logic_vector(31 downto 0);
    signal add_srcx_x1_at_entry_534 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1187_constant_part_of_offset : std_logic_vector(14 downto 0);
    signal array_obj_ref_1187_final_offset : std_logic_vector(14 downto 0);
    signal array_obj_ref_1187_offset_scale_factor_0 : std_logic_vector(14 downto 0);
    signal array_obj_ref_1187_offset_scale_factor_1 : std_logic_vector(14 downto 0);
    signal array_obj_ref_1187_offset_scale_factor_2 : std_logic_vector(14 downto 0);
    signal array_obj_ref_1187_resized_base_address : std_logic_vector(14 downto 0);
    signal array_obj_ref_1187_root_address : std_logic_vector(14 downto 0);
    signal array_obj_ref_1521_constant_part_of_offset : std_logic_vector(14 downto 0);
    signal array_obj_ref_1521_final_offset : std_logic_vector(14 downto 0);
    signal array_obj_ref_1521_offset_scale_factor_0 : std_logic_vector(14 downto 0);
    signal array_obj_ref_1521_offset_scale_factor_1 : std_logic_vector(14 downto 0);
    signal array_obj_ref_1521_offset_scale_factor_2 : std_logic_vector(14 downto 0);
    signal array_obj_ref_1521_resized_base_address : std_logic_vector(14 downto 0);
    signal array_obj_ref_1521_root_address : std_logic_vector(14 downto 0);
    signal array_obj_ref_283_constant_part_of_offset : std_logic_vector(14 downto 0);
    signal array_obj_ref_283_final_offset : std_logic_vector(14 downto 0);
    signal array_obj_ref_283_offset_scale_factor_0 : std_logic_vector(14 downto 0);
    signal array_obj_ref_283_offset_scale_factor_1 : std_logic_vector(14 downto 0);
    signal array_obj_ref_283_offset_scale_factor_2 : std_logic_vector(14 downto 0);
    signal array_obj_ref_283_resized_base_address : std_logic_vector(14 downto 0);
    signal array_obj_ref_283_root_address : std_logic_vector(14 downto 0);
    signal array_obj_ref_789_constant_part_of_offset : std_logic_vector(14 downto 0);
    signal array_obj_ref_789_final_offset : std_logic_vector(14 downto 0);
    signal array_obj_ref_789_offset_scale_factor_0 : std_logic_vector(14 downto 0);
    signal array_obj_ref_789_offset_scale_factor_1 : std_logic_vector(14 downto 0);
    signal array_obj_ref_789_offset_scale_factor_2 : std_logic_vector(14 downto 0);
    signal array_obj_ref_789_resized_base_address : std_logic_vector(14 downto 0);
    signal array_obj_ref_789_root_address : std_logic_vector(14 downto 0);
    signal arrayidx184_791 : std_logic_vector(31 downto 0);
    signal arrayidx250_1189 : std_logic_vector(31 downto 0);
    signal arrayidx375_1523 : std_logic_vector(31 downto 0);
    signal arrayidx_285 : std_logic_vector(31 downto 0);
    signal call100_373 : std_logic_vector(7 downto 0);
    signal call106_391 : std_logic_vector(7 downto 0);
    signal call10_85 : std_logic_vector(7 downto 0);
    signal call112_409 : std_logic_vector(7 downto 0);
    signal call120_445 : std_logic_vector(63 downto 0);
    signal call14_97 : std_logic_vector(7 downto 0);
    signal call19_110 : std_logic_vector(7 downto 0);
    signal call23_122 : std_logic_vector(7 downto 0);
    signal call28_136 : std_logic_vector(7 downto 0);
    signal call296_1345 : std_logic_vector(63 downto 0);
    signal call2_60 : std_logic_vector(7 downto 0);
    signal call32_148 : std_logic_vector(7 downto 0);
    signal call37_161 : std_logic_vector(7 downto 0);
    signal call41_173 : std_logic_vector(7 downto 0);
    signal call46_186 : std_logic_vector(7 downto 0);
    signal call5_72 : std_logic_vector(7 downto 0);
    signal call72_288 : std_logic_vector(7 downto 0);
    signal call76_301 : std_logic_vector(7 downto 0);
    signal call82_319 : std_logic_vector(7 downto 0);
    signal call88_337 : std_logic_vector(7 downto 0);
    signal call94_355 : std_logic_vector(7 downto 0);
    signal call_46 : std_logic_vector(7 downto 0);
    signal cmp158_650 : std_logic_vector(0 downto 0);
    signal cmp178_761 : std_logic_vector(0 downto 0);
    signal cmp196_864 : std_logic_vector(0 downto 0);
    signal cmp206_879 : std_logic_vector(0 downto 0);
    signal cmp217_925 : std_logic_vector(0 downto 0);
    signal cmp225_971 : std_logic_vector(0 downto 0);
    signal cmp245_1166 : std_logic_vector(0 downto 0);
    signal cmp261_1262 : std_logic_vector(0 downto 0);
    signal cmp274_1301 : std_logic_vector(0 downto 0);
    signal cmp284_1325 : std_logic_vector(0 downto 0);
    signal cmp369459_1460 : std_logic_vector(0 downto 0);
    signal cmp462_230 : std_logic_vector(0 downto 0);
    signal cond_1041 : std_logic_vector(31 downto 0);
    signal condx_xend_exec_guard_1000 : std_logic_vector(0 downto 0);
    signal condx_xend_exec_guard_933_delayed_1_0_1034 : std_logic_vector(0 downto 0);
    signal condx_xend_ifx_xend238_taken_1044 : std_logic_vector(0 downto 0);
    signal condx_xend_ifx_xend238_taken_949_delayed_10_0_1055 : std_logic_vector(0 downto 0);
    signal condx_xend_ifx_xend238_taken_997_delayed_1_0_1124 : std_logic_vector(0 downto 0);
    signal condx_xin_1031 : std_logic_vector(31 downto 0);
    signal conv102_377 : std_logic_vector(63 downto 0);
    signal conv108_395 : std_logic_vector(63 downto 0);
    signal conv114_413 : std_logic_vector(63 downto 0);
    signal conv11_89 : std_logic_vector(31 downto 0);
    signal conv121_1342 : std_logic_vector(63 downto 0);
    signal conv138_463 : std_logic_vector(31 downto 0);
    signal conv163_685 : std_logic_vector(31 downto 0);
    signal conv172445_742 : std_logic_vector(63 downto 0);
    signal conv17_101 : std_logic_vector(31 downto 0);
    signal conv193_855 : std_logic_vector(31 downto 0);
    signal conv1_51 : std_logic_vector(31 downto 0);
    signal conv20_114 : std_logic_vector(31 downto 0);
    signal conv210_916 : std_logic_vector(31 downto 0);
    signal conv221_953 : std_logic_vector(31 downto 0);
    signal conv257_1252 : std_logic_vector(31 downto 0);
    signal conv26_127 : std_logic_vector(15 downto 0);
    signal conv297_1350 : std_logic_vector(63 downto 0);
    signal conv29_140 : std_logic_vector(15 downto 0);
    signal conv305_1359 : std_logic_vector(7 downto 0);
    signal conv311_1369 : std_logic_vector(7 downto 0);
    signal conv317_1379 : std_logic_vector(7 downto 0);
    signal conv323_1389 : std_logic_vector(7 downto 0);
    signal conv329_1399 : std_logic_vector(7 downto 0);
    signal conv335_1409 : std_logic_vector(7 downto 0);
    signal conv341_1419 : std_logic_vector(7 downto 0);
    signal conv347_1429 : std_logic_vector(7 downto 0);
    signal conv35_152 : std_logic_vector(15 downto 0);
    signal conv380_1531 : std_logic_vector(7 downto 0);
    signal conv386_1541 : std_logic_vector(7 downto 0);
    signal conv38_165 : std_logic_vector(15 downto 0);
    signal conv392_1551 : std_logic_vector(7 downto 0);
    signal conv398_1561 : std_logic_vector(7 downto 0);
    signal conv3_64 : std_logic_vector(31 downto 0);
    signal conv404_1571 : std_logic_vector(7 downto 0);
    signal conv410_1581 : std_logic_vector(7 downto 0);
    signal conv416_1591 : std_logic_vector(7 downto 0);
    signal conv422_1601 : std_logic_vector(7 downto 0);
    signal conv44_177 : std_logic_vector(31 downto 0);
    signal conv47_190 : std_logic_vector(31 downto 0);
    signal conv61_209 : std_logic_vector(31 downto 0);
    signal conv63_213 : std_logic_vector(31 downto 0);
    signal conv73_292 : std_logic_vector(63 downto 0);
    signal conv78_305 : std_logic_vector(63 downto 0);
    signal conv84_323 : std_logic_vector(63 downto 0);
    signal conv8_76 : std_logic_vector(31 downto 0);
    signal conv90_341 : std_logic_vector(63 downto 0);
    signal conv96_359 : std_logic_vector(63 downto 0);
    signal exitcond7_1636 : std_logic_vector(0 downto 0);
    signal exitcond_433 : std_logic_vector(0 downto 0);
    signal iNsTr_16_488 : std_logic_vector(31 downto 0);
    signal iNsTr_28_1010_delayed_2_0_1142 : std_logic_vector(31 downto 0);
    signal iNsTr_28_600 : std_logic_vector(31 downto 0);
    signal iNsTr_28_at_entry_543 : std_logic_vector(31 downto 0);
    signal iNsTr_41_1272 : std_logic_vector(15 downto 0);
    signal ifx_xend186_exec_guard_660 : std_logic_vector(0 downto 0);
    signal ifx_xend186_ifx_xend238_taken_670 : std_logic_vector(0 downto 0);
    signal ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1047 : std_logic_vector(0 downto 0);
    signal ifx_xend238_exec_guard_1052 : std_logic_vector(0 downto 0);
    signal ifx_xend238_ifx_xend253_taken_1177 : std_logic_vector(0 downto 0);
    signal ifx_xend238_ifx_xthen247_taken_1171 : std_logic_vector(0 downto 0);
    signal ifx_xend253_whilex_xend_taken_1328 : std_logic_vector(0 downto 0);
    signal ifx_xend_exec_guard_673 : std_logic_vector(0 downto 0);
    signal ifx_xend_exec_guard_686_delayed_1_0_688 : std_logic_vector(0 downto 0);
    signal ifx_xend_exec_guard_693_delayed_1_0_698 : std_logic_vector(0 downto 0);
    signal ifx_xend_exec_guard_700_delayed_1_0_708 : std_logic_vector(0 downto 0);
    signal ifx_xend_exec_guard_705_delayed_2_0_716 : std_logic_vector(0 downto 0);
    signal ifx_xend_exec_guard_718_delayed_2_0_735 : std_logic_vector(0 downto 0);
    signal ifx_xend_exec_guard_725_delayed_2_0_745 : std_logic_vector(0 downto 0);
    signal ifx_xend_ifx_xthen180_taken_766 : std_logic_vector(0 downto 0);
    signal ifx_xend_ifx_xthen191_taken_772 : std_logic_vector(0 downto 0);
    signal ifx_xthen180_exec_guard_768_delayed_6_0_794 : std_logic_vector(0 downto 0);
    signal ifx_xthen180_exec_guard_775 : std_logic_vector(0 downto 0);
    signal ifx_xthen180_ifx_xthen191_taken_802 : std_logic_vector(0 downto 0);
    signal ifx_xthen180_ifx_xthen191_taken_807_delayed_12_0_835 : std_logic_vector(0 downto 0);
    signal ifx_xthen191_condx_xend_taken_896 : std_logic_vector(0 downto 0);
    signal ifx_xthen191_condx_xend_taken_911_delayed_1_0_993 : std_logic_vector(0 downto 0);
    signal ifx_xthen191_condx_xend_taken_918_delayed_2_0_1003 : std_logic_vector(0 downto 0);
    signal ifx_xthen191_exec_guard_807 : std_logic_vector(0 downto 0);
    signal ifx_xthen191_exec_guard_823_delayed_1_0_858 : std_logic_vector(0 downto 0);
    signal ifx_xthen191_exec_guard_829_delayed_1_0_867 : std_logic_vector(0 downto 0);
    signal ifx_xthen191_exec_guard_838_delayed_1_0_882 : std_logic_vector(0 downto 0);
    signal ifx_xthen191_exec_guard_845_delayed_1_0_891 : std_logic_vector(0 downto 0);
    signal ifx_xthen191_exec_guard_850_delayed_1_0_899 : std_logic_vector(0 downto 0);
    signal ifx_xthen191_landx_xlhsx_xtrue208_taken_905 : std_logic_vector(0 downto 0);
    signal ifx_xthen247_exec_guard_1180 : std_logic_vector(0 downto 0);
    signal ifx_xthen247_ifx_xend253_taken_1207 : std_logic_vector(0 downto 0);
    signal inc162_680 : std_logic_vector(7 downto 0);
    signal inc240_1149 : std_logic_vector(31 downto 0);
    signal inc242_1159 : std_logic_vector(7 downto 0);
    signal inc252_1204 : std_logic_vector(31 downto 0);
    signal inc265_1139_delayed_1_0_1289 : std_logic_vector(15 downto 0);
    signal inc265_1268 : std_logic_vector(15 downto 0);
    signal inc268_1278 : std_logic_vector(15 downto 0);
    signal inc278_1305 : std_logic_vector(15 downto 0);
    signal inc278x_xo0x_x1_1313 : std_logic_vector(15 downto 0);
    signal inc442_1631 : std_logic_vector(31 downto 0);
    signal inc_428 : std_logic_vector(31 downto 0);
    signal input_byte_countx_x1_615 : std_logic_vector(7 downto 0);
    signal input_byte_countx_x1_at_entry_558 : std_logic_vector(7 downto 0);
    signal input_byte_countx_x2454_1088 : std_logic_vector(7 downto 0);
    signal input_byte_countx_x2x_xph_832 : std_logic_vector(7 downto 0);
    signal input_wordx_x0456_1070 : std_logic_vector(63 downto 0);
    signal input_wordx_x0x_xph_850 : std_logic_vector(63 downto 0);
    signal input_wordx_x1_640 : std_logic_vector(63 downto 0);
    signal input_wordx_x1_707_delayed_2_0_719 : std_logic_vector(63 downto 0);
    signal input_wordx_x1_at_entry_583 : std_logic_vector(63 downto 0);
    signal input_wordx_x1_at_entry_583_644_buffered : std_logic_vector(63 downto 0);
    signal ix_x0463_269 : std_logic_vector(31 downto 0);
    signal ix_x1460_1507 : std_logic_vector(31 downto 0);
    signal landx_xlhsx_xtrue208_condx_xend_taken_921_delayed_1_0_1010 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue208_condx_xend_taken_942 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue208_exec_guard_863_delayed_1_0_919 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_928 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_936 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue208_exec_guard_908 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue208_landx_xlhsx_xtrue219_taken_933 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue219_condx_xend_taken_924_delayed_1_0_1017 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue219_condx_xend_taken_990 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue219_exec_guard_894_delayed_1_0_965 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue219_exec_guard_900_delayed_1_0_974 : std_logic_vector(0 downto 0);
    signal landx_xlhsx_xtrue219_exec_guard_945 : std_logic_vector(0 downto 0);
    signal mul143_468 : std_logic_vector(31 downto 0);
    signal mul145_478 : std_logic_vector(31 downto 0);
    signal mul164_695 : std_logic_vector(31 downto 0);
    signal mul230_526 : std_logic_vector(31 downto 0);
    signal mul233_531 : std_logic_vector(31 downto 0);
    signal mul58_205 : std_logic_vector(31 downto 0);
    signal mul64_218 : std_logic_vector(31 downto 0);
    signal mul67_223 : std_logic_vector(31 downto 0);
    signal mul_200 : std_logic_vector(31 downto 0);
    signal o0x_x1_1155_delayed_3_0_1308 : std_logic_vector(15 downto 0);
    signal o0x_x1_620 : std_logic_vector(15 downto 0);
    signal o0x_x1_at_entry_563 : std_logic_vector(15 downto 0);
    signal o1x_x0_1286 : std_logic_vector(15 downto 0);
    signal o1x_x1_1134_delayed_2_0_1281 : std_logic_vector(15 downto 0);
    signal o1x_x1_625 : std_logic_vector(15 downto 0);
    signal o1x_x1_860_delayed_1_0_911 : std_logic_vector(15 downto 0);
    signal o1x_x1_at_entry_568 : std_logic_vector(15 downto 0);
    signal o1x_x2_1320 : std_logic_vector(15 downto 0);
    signal o2x_x0_1296 : std_logic_vector(15 downto 0);
    signal o2x_x1_630 : std_logic_vector(15 downto 0);
    signal o2x_x1_885_delayed_2_0_948 : std_logic_vector(15 downto 0);
    signal o2x_x1_at_entry_573 : std_logic_vector(15 downto 0);
    signal orx_xcond_888 : std_logic_vector(0 downto 0);
    signal output_byte_countx_x0_1017_delayed_2_0_1152 : std_logic_vector(7 downto 0);
    signal output_byte_countx_x0_610 : std_logic_vector(7 downto 0);
    signal output_byte_countx_x0_at_entry_553 : std_logic_vector(7 downto 0);
    signal output_byte_countx_x1_1235 : std_logic_vector(7 downto 0);
    signal ptr_deref_1192_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1192_resized_base_address : std_logic_vector(14 downto 0);
    signal ptr_deref_1192_root_address : std_logic_vector(14 downto 0);
    signal ptr_deref_1192_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1192_word_address_0 : std_logic_vector(14 downto 0);
    signal ptr_deref_1192_word_offset_0 : std_logic_vector(14 downto 0);
    signal ptr_deref_1526_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1526_resized_base_address : std_logic_vector(14 downto 0);
    signal ptr_deref_1526_root_address : std_logic_vector(14 downto 0);
    signal ptr_deref_1526_word_address_0 : std_logic_vector(14 downto 0);
    signal ptr_deref_1526_word_offset_0 : std_logic_vector(14 downto 0);
    signal ptr_deref_420_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_420_resized_base_address : std_logic_vector(14 downto 0);
    signal ptr_deref_420_root_address : std_logic_vector(14 downto 0);
    signal ptr_deref_420_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_420_word_address_0 : std_logic_vector(14 downto 0);
    signal ptr_deref_420_word_offset_0 : std_logic_vector(14 downto 0);
    signal ptr_deref_491_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_491_resized_base_address : std_logic_vector(14 downto 0);
    signal ptr_deref_491_root_address : std_logic_vector(14 downto 0);
    signal ptr_deref_491_word_address_0 : std_logic_vector(14 downto 0);
    signal ptr_deref_491_word_offset_0 : std_logic_vector(14 downto 0);
    signal ptr_deref_798_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_798_resized_base_address : std_logic_vector(14 downto 0);
    signal ptr_deref_798_root_address : std_logic_vector(14 downto 0);
    signal ptr_deref_798_word_address_0 : std_logic_vector(14 downto 0);
    signal ptr_deref_798_word_offset_0 : std_logic_vector(14 downto 0);
    signal sh_prom_713 : std_logic_vector(63 downto 0);
    signal shl105_388 : std_logic_vector(63 downto 0);
    signal shl111_406 : std_logic_vector(63 downto 0);
    signal shl169_728_delayed_2_0_748 : std_logic_vector(63 downto 0);
    signal shl169_732 : std_logic_vector(63 downto 0);
    signal shl175_667 : std_logic_vector(63 downto 0);
    signal shl18_107 : std_logic_vector(31 downto 0);
    signal shl27_133 : std_logic_vector(15 downto 0);
    signal shl36_158 : std_logic_vector(15 downto 0);
    signal shl45_183 : std_logic_vector(31 downto 0);
    signal shl75_298 : std_logic_vector(63 downto 0);
    signal shl81_316 : std_logic_vector(63 downto 0);
    signal shl87_334 : std_logic_vector(63 downto 0);
    signal shl93_352 : std_logic_vector(63 downto 0);
    signal shl99_370 : std_logic_vector(63 downto 0);
    signal shl9_82 : std_logic_vector(31 downto 0);
    signal shl_57 : std_logic_vector(31 downto 0);
    signal shr130444_457 : std_logic_vector(31 downto 0);
    signal shr166_725 : std_logic_vector(63 downto 0);
    signal shr308_1365 : std_logic_vector(63 downto 0);
    signal shr314_1375 : std_logic_vector(63 downto 0);
    signal shr320_1385 : std_logic_vector(63 downto 0);
    signal shr326_1395 : std_logic_vector(63 downto 0);
    signal shr332_1405 : std_logic_vector(63 downto 0);
    signal shr338_1415 : std_logic_vector(63 downto 0);
    signal shr344_1425 : std_logic_vector(63 downto 0);
    signal shr383_1537 : std_logic_vector(63 downto 0);
    signal shr389_1547 : std_logic_vector(63 downto 0);
    signal shr395_1557 : std_logic_vector(63 downto 0);
    signal shr401_1567 : std_logic_vector(63 downto 0);
    signal shr407_1577 : std_logic_vector(63 downto 0);
    signal shr413_1587 : std_logic_vector(63 downto 0);
    signal shr419_1597 : std_logic_vector(63 downto 0);
    signal sub165_705 : std_logic_vector(31 downto 0);
    signal sub204_498 : std_logic_vector(31 downto 0);
    signal sub205_503 : std_logic_vector(31 downto 0);
    signal sub215_509 : std_logic_vector(31 downto 0);
    signal sub216_514 : std_logic_vector(31 downto 0);
    signal sub224_520 : std_logic_vector(31 downto 0);
    signal sub301_1355 : std_logic_vector(63 downto 0);
    signal sub_451 : std_logic_vector(31 downto 0);
    signal target_out_offsetx_x0_1139 : std_logic_vector(31 downto 0);
    signal target_out_offsetx_x1_595 : std_logic_vector(31 downto 0);
    signal target_out_offsetx_x1_890_delayed_2_0_956 : std_logic_vector(31 downto 0);
    signal target_out_offsetx_x1_904_delayed_3_0_980 : std_logic_vector(31 downto 0);
    signal target_out_offsetx_x1_at_entry_539 : std_logic_vector(31 downto 0);
    signal target_out_offsetx_x1_at_entry_539_599_buffered : std_logic_vector(31 downto 0);
    signal tmp10_253 : std_logic_vector(31 downto 0);
    signal tmp11_259 : std_logic_vector(0 downto 0);
    signal tmp155_492 : std_logic_vector(63 downto 0);
    signal tmp185_799 : std_logic_vector(63 downto 0);
    signal tmp1_1476 : std_logic_vector(31 downto 0);
    signal tmp2_1480 : std_logic_vector(31 downto 0);
    signal tmp376_1527 : std_logic_vector(63 downto 0);
    signal tmp3_1485 : std_logic_vector(31 downto 0);
    signal tmp4_1491 : std_logic_vector(31 downto 0);
    signal tmp5_1497 : std_logic_vector(0 downto 0);
    signal tmp8_242 : std_logic_vector(31 downto 0);
    signal tmp9_247 : std_logic_vector(31 downto 0);
    signal tmp_1471 : std_logic_vector(31 downto 0);
    signal type_cast_1025_wire : std_logic_vector(31 downto 0);
    signal type_cast_1027_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1039_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1059_wire : std_logic_vector(63 downto 0);
    signal type_cast_105_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1061_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1067_wire : std_logic_vector(63 downto 0);
    signal type_cast_1073_1073_delayed_2_0_1211 : std_logic_vector(31 downto 0);
    signal type_cast_1078_wire : std_logic_vector(7 downto 0);
    signal type_cast_1080_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1096_wire : std_logic_vector(31 downto 0);
    signal type_cast_1098_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1110_wire : std_logic_vector(63 downto 0);
    signal type_cast_1112_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1113_1113_delayed_2_0_1256 : std_logic_vector(31 downto 0);
    signal type_cast_1118_wire : std_logic_vector(63 downto 0);
    signal type_cast_1128_wire : std_logic_vector(31 downto 0);
    signal type_cast_1130_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1136_wire : std_logic_vector(31 downto 0);
    signal type_cast_1147_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1157_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1164_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1202_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1215_wire : std_logic_vector(31 downto 0);
    signal type_cast_1219_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1227_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1230_wire : std_logic_vector(7 downto 0);
    signal type_cast_1232_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1240_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1243_wire : std_logic_vector(63 downto 0);
    signal type_cast_1245_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1259_wire : std_logic_vector(31 downto 0);
    signal type_cast_1266_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1276_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1294_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1317_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_131_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1340_wire : std_logic_vector(63 downto 0);
    signal type_cast_1348_wire : std_logic_vector(63 downto 0);
    signal type_cast_1363_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1373_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1383_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1393_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1403_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1413_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1423_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1458_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1489_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1495_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1502_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1511_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1513_wire : std_logic_vector(31 downto 0);
    signal type_cast_1535_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1545_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1555_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1565_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_156_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1575_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1585_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1595_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1629_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_181_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_227_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_251_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_257_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_264_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_273_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_275_wire : std_logic_vector(31 downto 0);
    signal type_cast_296_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_314_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_332_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_350_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_368_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_386_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_404_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_426_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_455_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_461_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_496_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_507_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_518_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_524_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_542_wire : std_logic_vector(31 downto 0);
    signal type_cast_55_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_586_wire : std_logic_vector(63 downto 0);
    signal type_cast_593_wire : std_logic_vector(31 downto 0);
    signal type_cast_598_wire : std_logic_vector(31 downto 0);
    signal type_cast_603_wire : std_logic_vector(31 downto 0);
    signal type_cast_608_wire : std_logic_vector(31 downto 0);
    signal type_cast_613_wire : std_logic_vector(7 downto 0);
    signal type_cast_618_wire : std_logic_vector(7 downto 0);
    signal type_cast_623_wire : std_logic_vector(15 downto 0);
    signal type_cast_628_wire : std_logic_vector(15 downto 0);
    signal type_cast_633_wire : std_logic_vector(15 downto 0);
    signal type_cast_638_wire : std_logic_vector(63 downto 0);
    signal type_cast_643_wire : std_logic_vector(63 downto 0);
    signal type_cast_665_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_678_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_693_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_702_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_730_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_740_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_759_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_780_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_80_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_811_wire : std_logic_vector(31 downto 0);
    signal type_cast_814_wire : std_logic_vector(31 downto 0);
    signal type_cast_816_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_824_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_827_wire : std_logic_vector(7 downto 0);
    signal type_cast_829_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_835_835_delayed_1_0_872 : std_logic_vector(31 downto 0);
    signal type_cast_839_wire : std_logic_vector(63 downto 0);
    signal type_cast_841_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_847_wire : std_logic_vector(63 downto 0);
    signal type_cast_876_wire : std_logic_vector(31 downto 0);
    signal type_cast_920_920_delayed_3_0_1007 : std_logic_vector(31 downto 0);
    signal type_cast_923_923_delayed_3_0_1014 : std_logic_vector(31 downto 0);
    signal type_cast_963_963_delayed_2_0_1074 : std_logic_vector(7 downto 0);
    signal type_cast_975_975_delayed_2_0_1092 : std_logic_vector(31 downto 0);
    signal umax6_1504 : std_logic_vector(31 downto 0);
    signal umax_266 : std_logic_vector(31 downto 0);
    signal valuex_x0448450_1121 : std_logic_vector(63 downto 0);
    signal valuex_x1_635 : std_logic_vector(63 downto 0);
    signal valuex_x1_at_entry_578 : std_logic_vector(63 downto 0);
    signal valuex_x2_1248 : std_logic_vector(63 downto 0);
    signal whilex_xbody_ifx_xend186_taken_657 : std_logic_vector(0 downto 0);
    signal whilex_xbody_ifx_xend_taken_653 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    add_outx_x1_at_entry_548 <= "00000000000000000000000000000000";
    add_srcx_x1_at_entry_534 <= "00000000000000000000000000000000";
    array_obj_ref_1187_constant_part_of_offset <= "100000000000000";
    array_obj_ref_1187_offset_scale_factor_0 <= "100000000000000";
    array_obj_ref_1187_offset_scale_factor_1 <= "100000000000000";
    array_obj_ref_1187_offset_scale_factor_2 <= "000000000000001";
    array_obj_ref_1187_resized_base_address <= "000000000000000";
    array_obj_ref_1521_constant_part_of_offset <= "100000000000000";
    array_obj_ref_1521_offset_scale_factor_0 <= "100000000000000";
    array_obj_ref_1521_offset_scale_factor_1 <= "100000000000000";
    array_obj_ref_1521_offset_scale_factor_2 <= "000000000000001";
    array_obj_ref_1521_resized_base_address <= "000000000000000";
    array_obj_ref_283_constant_part_of_offset <= "000000000000000";
    array_obj_ref_283_offset_scale_factor_0 <= "100000000000000";
    array_obj_ref_283_offset_scale_factor_1 <= "100000000000000";
    array_obj_ref_283_offset_scale_factor_2 <= "000000000000001";
    array_obj_ref_283_resized_base_address <= "000000000000000";
    array_obj_ref_789_constant_part_of_offset <= "000000000000000";
    array_obj_ref_789_offset_scale_factor_0 <= "100000000000000";
    array_obj_ref_789_offset_scale_factor_1 <= "100000000000000";
    array_obj_ref_789_offset_scale_factor_2 <= "000000000000001";
    array_obj_ref_789_resized_base_address <= "000000000000000";
    iNsTr_16_488 <= "00000000000000000000000000000000";
    iNsTr_28_at_entry_543 <= "00000000000000000000000000000000";
    input_byte_countx_x1_at_entry_558 <= "00000000";
    o0x_x1_at_entry_563 <= "0000000000000000";
    o1x_x1_at_entry_568 <= "0000000000000000";
    o2x_x1_at_entry_573 <= "0000000000000000";
    output_byte_countx_x0_at_entry_553 <= "00000000";
    ptr_deref_1192_word_offset_0 <= "000000000000000";
    ptr_deref_1526_word_offset_0 <= "000000000000000";
    ptr_deref_420_word_offset_0 <= "000000000000000";
    ptr_deref_491_word_offset_0 <= "000000000000000";
    ptr_deref_798_word_offset_0 <= "000000000000000";
    type_cast_1027_wire_constant <= "00000000000000000000000000000000";
    type_cast_1039_wire_constant <= "00000000000000000000000000000001";
    type_cast_105_wire_constant <= "00000000000000000000000000001000";
    type_cast_1061_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1080_wire_constant <= "00000000";
    type_cast_1098_wire_constant <= "00000000000000000000000000000000";
    type_cast_1112_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1130_wire_constant <= "00000000000000000000000000000000";
    type_cast_1147_wire_constant <= "00000000000000000000000000000001";
    type_cast_1157_wire_constant <= "00000001";
    type_cast_1164_wire_constant <= "00001000";
    type_cast_1202_wire_constant <= "00000000000000000000000000000001";
    type_cast_1219_wire_constant <= "00000000000000000000000000000000";
    type_cast_1227_wire_constant <= "00000000";
    type_cast_1232_wire_constant <= "00000000";
    type_cast_1240_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1245_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1266_wire_constant <= "0000000000000001";
    type_cast_1276_wire_constant <= "0000000000000001";
    type_cast_1294_wire_constant <= "0000000000000000";
    type_cast_1317_wire_constant <= "0000000000000000";
    type_cast_131_wire_constant <= "0000000000001000";
    type_cast_1363_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1373_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1383_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1393_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1403_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1413_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1423_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1458_wire_constant <= "00000000000000000000000000000111";
    type_cast_1489_wire_constant <= "00000000000000000000000000000011";
    type_cast_1495_wire_constant <= "00000000000000000000000000000001";
    type_cast_1502_wire_constant <= "00000000000000000000000000000001";
    type_cast_1511_wire_constant <= "00000000000000000000000000000000";
    type_cast_1535_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1545_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1555_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1565_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_156_wire_constant <= "0000000000001000";
    type_cast_1575_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1585_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1595_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1629_wire_constant <= "00000000000000000000000000000001";
    type_cast_181_wire_constant <= "00000000000000000000000000001000";
    type_cast_227_wire_constant <= "00000000000000000000000000000111";
    type_cast_251_wire_constant <= "00000000000000000000000000000011";
    type_cast_257_wire_constant <= "00000000000000000000000000000001";
    type_cast_264_wire_constant <= "00000000000000000000000000000001";
    type_cast_273_wire_constant <= "00000000000000000000000000000000";
    type_cast_296_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_314_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_332_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_350_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_368_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_386_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_404_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_426_wire_constant <= "00000000000000000000000000000001";
    type_cast_455_wire_constant <= "00000000000000000000000000000001";
    type_cast_461_wire_constant <= "00000000000000000000000011111111";
    type_cast_496_wire_constant <= "11111111111111111111111111111111";
    type_cast_507_wire_constant <= "11111111111111111111111111111111";
    type_cast_518_wire_constant <= "11111111111111111111111111111111";
    type_cast_524_wire_constant <= "00000000000000000000000111111110";
    type_cast_55_wire_constant <= "00000000000000000000000000001000";
    type_cast_665_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_678_wire_constant <= "00000001";
    type_cast_693_wire_constant <= "00000000000000000000000000000011";
    type_cast_702_wire_constant <= "00000000000000000000000000111000";
    type_cast_730_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_740_wire_constant <= "0000000000000000000000000000000000000000000000000000000011111111";
    type_cast_759_wire_constant <= "00001000";
    type_cast_780_wire_constant <= "00000000000000000000000000000001";
    type_cast_80_wire_constant <= "00000000000000000000000000001000";
    type_cast_816_wire_constant <= "00000000000000000000000000000000";
    type_cast_824_wire_constant <= "00000000";
    type_cast_829_wire_constant <= "00000000";
    type_cast_841_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    valuex_x1_at_entry_578 <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_1507: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1511_wire_constant & type_cast_1513_wire;
      req <= phi_stmt_1507_req_0 & phi_stmt_1507_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1507",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1507_ack_0,
          idata => idata,
          odata => ix_x1460_1507,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1507
    phi_stmt_269: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_273_wire_constant & type_cast_275_wire;
      req <= phi_stmt_269_req_0 & phi_stmt_269_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_269",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_269_ack_0,
          idata => idata,
          odata => ix_x0463_269,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_269
    phi_stmt_539: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_542_wire;
      req(0) <= phi_stmt_539_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_539",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_539_ack_0,
          idata => idata,
          odata => target_out_offsetx_x1_at_entry_539,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_539
    phi_stmt_583: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_586_wire;
      req(0) <= phi_stmt_583_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_583",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_583_ack_0,
          idata => idata,
          odata => input_wordx_x1_at_entry_583,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_583
    phi_stmt_590: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_593_wire & add_srcx_x1_at_entry_534;
      req <= phi_stmt_590_req_0 & phi_stmt_590_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_590",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_590_ack_0,
          idata => idata,
          odata => add_srcx_x1_590,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_590
    phi_stmt_595: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_598_wire & target_out_offsetx_x1_at_entry_539_599_buffered;
      req <= phi_stmt_595_req_0 & phi_stmt_595_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_595",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_595_ack_0,
          idata => idata,
          odata => target_out_offsetx_x1_595,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_595
    phi_stmt_600: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_603_wire & iNsTr_28_at_entry_543;
      req <= phi_stmt_600_req_0 & phi_stmt_600_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_600",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_600_ack_0,
          idata => idata,
          odata => iNsTr_28_600,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_600
    phi_stmt_605: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_608_wire & add_outx_x1_at_entry_548;
      req <= phi_stmt_605_req_0 & phi_stmt_605_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_605",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_605_ack_0,
          idata => idata,
          odata => add_outx_x1_605,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_605
    phi_stmt_610: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_613_wire & output_byte_countx_x0_at_entry_553;
      req <= phi_stmt_610_req_0 & phi_stmt_610_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_610",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_610_ack_0,
          idata => idata,
          odata => output_byte_countx_x0_610,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_610
    phi_stmt_615: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_618_wire & input_byte_countx_x1_at_entry_558;
      req <= phi_stmt_615_req_0 & phi_stmt_615_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_615",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_615_ack_0,
          idata => idata,
          odata => input_byte_countx_x1_615,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_615
    phi_stmt_620: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_623_wire & o0x_x1_at_entry_563;
      req <= phi_stmt_620_req_0 & phi_stmt_620_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_620",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_620_ack_0,
          idata => idata,
          odata => o0x_x1_620,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_620
    phi_stmt_625: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_628_wire & o1x_x1_at_entry_568;
      req <= phi_stmt_625_req_0 & phi_stmt_625_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_625",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_625_ack_0,
          idata => idata,
          odata => o1x_x1_625,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_625
    phi_stmt_630: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_633_wire & o2x_x1_at_entry_573;
      req <= phi_stmt_630_req_0 & phi_stmt_630_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_630",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_630_ack_0,
          idata => idata,
          odata => o2x_x1_630,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_630
    phi_stmt_635: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_638_wire & valuex_x1_at_entry_578;
      req <= phi_stmt_635_req_0 & phi_stmt_635_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_635",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_635_ack_0,
          idata => idata,
          odata => valuex_x1_635,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_635
    phi_stmt_640: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_643_wire & input_wordx_x1_at_entry_583_644_buffered;
      req <= phi_stmt_640_req_0 & phi_stmt_640_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_640",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_640_ack_0,
          idata => idata,
          odata => input_wordx_x1_640,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_640
    -- flow-through select operator MUX_1028_inst
    MUX_1028_wire <= type_cast_1025_wire when (landx_xlhsx_xtrue219_condx_xend_taken_924_delayed_1_0_1017(0) /=  '0') else type_cast_1027_wire_constant;
    -- flow-through select operator MUX_1029_inst
    MUX_1029_wire <= type_cast_923_923_delayed_3_0_1014 when (landx_xlhsx_xtrue208_condx_xend_taken_921_delayed_1_0_1010(0) /=  '0') else MUX_1028_wire;
    -- flow-through select operator MUX_1030_inst
    condx_xin_1031 <= type_cast_920_920_delayed_3_0_1007 when (ifx_xthen191_condx_xend_taken_918_delayed_2_0_1003(0) /=  '0') else MUX_1029_wire;
    MUX_1062_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1062_inst_req_0;
      MUX_1062_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1062_inst_req_1;
      MUX_1062_inst_ack_1<= update_ack(0);
      MUX_1062_inst: SelectSplitProtocol generic map(name => "MUX_1062_inst", data_width => 64, buffering => 12, flow_through => false, full_rate => true) -- 
        port map( x => type_cast_1059_wire, y => type_cast_1061_wire_constant, sel => ifx_xend186_ifx_xend238_taken_670, z => MUX_957_957_delayed_12_0_1063, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_1069_inst
    input_wordx_x0456_1070 <= type_cast_1067_wire when (condx_xend_ifx_xend238_taken_949_delayed_10_0_1055(0) /=  '0') else MUX_957_957_delayed_12_0_1063;
    MUX_1081_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1081_inst_req_0;
      MUX_1081_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1081_inst_req_1;
      MUX_1081_inst_ack_1<= update_ack(0);
      MUX_1081_inst: SelectSplitProtocol generic map(name => "MUX_1081_inst", data_width => 8, buffering => 2, flow_through => false, full_rate => true) -- 
        port map( x => type_cast_1078_wire, y => type_cast_1080_wire_constant, sel => ifx_xend186_ifx_xend238_taken_670, z => MUX_969_969_delayed_2_0_1082, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_1087_inst
    input_byte_countx_x2454_1088 <= type_cast_963_963_delayed_2_0_1074 when (condx_xend_ifx_xend238_taken_1044(0) /=  '0') else MUX_969_969_delayed_2_0_1082;
    MUX_1099_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1099_inst_req_0;
      MUX_1099_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1099_inst_req_1;
      MUX_1099_inst_ack_1<= update_ack(0);
      MUX_1099_inst: SelectSplitProtocol generic map(name => "MUX_1099_inst", data_width => 32, buffering => 2, flow_through => false, full_rate => true) -- 
        port map( x => type_cast_1096_wire, y => type_cast_1098_wire_constant, sel => ifx_xend186_ifx_xend238_taken_670, z => MUX_981_981_delayed_2_0_1100, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_1105_inst
    add_srcx_x0452_1106 <= type_cast_975_975_delayed_2_0_1092 when (condx_xend_ifx_xend238_taken_1044(0) /=  '0') else MUX_981_981_delayed_2_0_1100;
    MUX_1113_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1113_inst_req_0;
      MUX_1113_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1113_inst_req_1;
      MUX_1113_inst_ack_1<= update_ack(0);
      MUX_1113_inst: SelectSplitProtocol generic map(name => "MUX_1113_inst", data_width => 64, buffering => 2, flow_through => false, full_rate => true) -- 
        port map( x => type_cast_1110_wire, y => type_cast_1112_wire_constant, sel => ifx_xend186_ifx_xend238_taken_670, z => MUX_993_993_delayed_2_0_1114, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_1120_inst
    valuex_x0448450_1121 <= type_cast_1118_wire when (condx_xend_ifx_xend238_taken_1044(0) /=  '0') else MUX_993_993_delayed_2_0_1114;
    MUX_1131_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_1131_inst_req_0;
      MUX_1131_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_1131_inst_req_1;
      MUX_1131_inst_ack_1<= update_ack(0);
      MUX_1131_inst: SelectSplitProtocol generic map(name => "MUX_1131_inst", data_width => 32, buffering => 3, flow_through => false, full_rate => true) -- 
        port map( x => type_cast_1128_wire, y => type_cast_1130_wire_constant, sel => ifx_xend186_ifx_xend238_taken_670, z => MUX_1005_1005_delayed_3_0_1132, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_1138_inst
    target_out_offsetx_x0_1139 <= type_cast_1136_wire when (condx_xend_ifx_xend238_taken_997_delayed_1_0_1124(0) /=  '0') else MUX_1005_1005_delayed_3_0_1132;
    -- flow-through select operator MUX_1220_inst
    MUX_1220_wire <= type_cast_1073_1073_delayed_2_0_1211 when (ifx_xend238_ifx_xend253_taken_1177(0) /=  '0') else type_cast_1219_wire_constant;
    -- flow-through select operator MUX_1221_inst
    add_outx_x0_1222 <= type_cast_1215_wire when (ifx_xthen247_ifx_xend253_taken_1207(0) /=  '0') else MUX_1220_wire;
    -- flow-through select operator MUX_1233_inst
    MUX_1233_wire <= type_cast_1230_wire when (ifx_xend238_ifx_xend253_taken_1177(0) /=  '0') else type_cast_1232_wire_constant;
    -- flow-through select operator MUX_1234_inst
    output_byte_countx_x1_1235 <= type_cast_1227_wire_constant when (ifx_xthen247_ifx_xend253_taken_1207(0) /=  '0') else MUX_1233_wire;
    -- flow-through select operator MUX_1246_inst
    MUX_1246_wire <= type_cast_1243_wire when (ifx_xend238_ifx_xend253_taken_1177(0) /=  '0') else type_cast_1245_wire_constant;
    -- flow-through select operator MUX_1247_inst
    valuex_x2_1248 <= type_cast_1240_wire_constant when (ifx_xthen247_ifx_xend253_taken_1207(0) /=  '0') else MUX_1246_wire;
    -- flow-through select operator MUX_1295_inst
    o2x_x0_1296 <= inc265_1139_delayed_1_0_1289 when (cmp261_1262(0) /=  '0') else type_cast_1294_wire_constant;
    -- flow-through select operator MUX_1319_inst
    o1x_x2_1320 <= type_cast_1317_wire_constant when (cmp274_1301(0) /=  '0') else o1x_x0_1286;
    -- flow-through select operator MUX_1503_inst
    umax6_1504 <= tmp4_1491 when (tmp5_1497(0) /=  '0') else type_cast_1502_wire_constant;
    -- flow-through select operator MUX_265_inst
    umax_266 <= tmp10_253 when (tmp11_259(0) /=  '0') else type_cast_264_wire_constant;
    -- flow-through select operator MUX_817_inst
    MUX_817_wire <= type_cast_814_wire when (ifx_xend_ifx_xthen191_taken_772(0) /=  '0') else type_cast_816_wire_constant;
    -- flow-through select operator MUX_818_inst
    add_srcx_x0x_xph_819 <= type_cast_811_wire when (ifx_xthen180_ifx_xthen191_taken_802(0) /=  '0') else MUX_817_wire;
    -- flow-through select operator MUX_830_inst
    MUX_830_wire <= type_cast_827_wire when (ifx_xend_ifx_xthen191_taken_772(0) /=  '0') else type_cast_829_wire_constant;
    -- flow-through select operator MUX_831_inst
    input_byte_countx_x2x_xph_832 <= type_cast_824_wire_constant when (ifx_xthen180_ifx_xthen191_taken_802(0) /=  '0') else MUX_830_wire;
    MUX_842_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_842_inst_req_0;
      MUX_842_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_842_inst_req_1;
      MUX_842_inst_ack_1<= update_ack(0);
      MUX_842_inst: SelectSplitProtocol generic map(name => "MUX_842_inst", data_width => 64, buffering => 12, flow_through => false, full_rate => true) -- 
        port map( x => type_cast_839_wire, y => type_cast_841_wire_constant, sel => ifx_xend_ifx_xthen191_taken_772, z => MUX_815_815_delayed_12_0_843, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_849_inst
    input_wordx_x0x_xph_850 <= type_cast_847_wire when (ifx_xthen180_ifx_xthen191_taken_807_delayed_12_0_835(0) /=  '0') else MUX_815_815_delayed_12_0_843;
    -- flow-through select operator MUX_986_inst
    add234x_xtarget_out_offsetx_x1_987 <= add234_903_delayed_1_0_977 when (cmp225_971(0) /=  '0') else target_out_offsetx_x1_904_delayed_3_0_980;
    W_add234_903_delayed_1_0_975_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add234_903_delayed_1_0_975_inst_req_0;
      W_add234_903_delayed_1_0_975_inst_ack_0<= wack(0);
      rreq(0) <= W_add234_903_delayed_1_0_975_inst_req_1;
      W_add234_903_delayed_1_0_975_inst_ack_1<= rack(0);
      W_add234_903_delayed_1_0_975_inst : InterlockBuffer generic map ( -- 
        name => "W_add234_903_delayed_1_0_975_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add234_962,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add234_903_delayed_1_0_977,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add_outx_x1_1059_delayed_2_0_1195_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_outx_x1_1059_delayed_2_0_1195_inst_req_0;
      W_add_outx_x1_1059_delayed_2_0_1195_inst_ack_0<= wack(0);
      rreq(0) <= W_add_outx_x1_1059_delayed_2_0_1195_inst_req_1;
      W_add_outx_x1_1059_delayed_2_0_1195_inst_ack_1<= rack(0);
      W_add_outx_x1_1059_delayed_2_0_1195_inst : InterlockBuffer generic map ( -- 
        name => "W_add_outx_x1_1059_delayed_2_0_1195_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x1_605,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_outx_x1_1059_delayed_2_0_1197,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_condx_xend_exec_guard_933_delayed_1_0_1032_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_condx_xend_exec_guard_933_delayed_1_0_1032_inst_req_0;
      W_condx_xend_exec_guard_933_delayed_1_0_1032_inst_ack_0<= wack(0);
      rreq(0) <= W_condx_xend_exec_guard_933_delayed_1_0_1032_inst_req_1;
      W_condx_xend_exec_guard_933_delayed_1_0_1032_inst_ack_1<= rack(0);
      W_condx_xend_exec_guard_933_delayed_1_0_1032_inst : InterlockBuffer generic map ( -- 
        name => "W_condx_xend_exec_guard_933_delayed_1_0_1032_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => condx_xend_exec_guard_1000,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => condx_xend_exec_guard_933_delayed_1_0_1034,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_condx_xend_ifx_xend238_taken_1042_inst
    process(condx_xend_exec_guard_1000) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := condx_xend_exec_guard_1000(0 downto 0);
      condx_xend_ifx_xend238_taken_1044 <= tmp_var; -- 
    end process;
    W_condx_xend_ifx_xend238_taken_949_delayed_10_0_1053_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_condx_xend_ifx_xend238_taken_949_delayed_10_0_1053_inst_req_0;
      W_condx_xend_ifx_xend238_taken_949_delayed_10_0_1053_inst_ack_0<= wack(0);
      rreq(0) <= W_condx_xend_ifx_xend238_taken_949_delayed_10_0_1053_inst_req_1;
      W_condx_xend_ifx_xend238_taken_949_delayed_10_0_1053_inst_ack_1<= rack(0);
      W_condx_xend_ifx_xend238_taken_949_delayed_10_0_1053_inst : InterlockBuffer generic map ( -- 
        name => "W_condx_xend_ifx_xend238_taken_949_delayed_10_0_1053_inst",
        buffer_size => 10,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => condx_xend_ifx_xend238_taken_1044,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => condx_xend_ifx_xend238_taken_949_delayed_10_0_1055,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_condx_xend_ifx_xend238_taken_997_delayed_1_0_1122_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_condx_xend_ifx_xend238_taken_997_delayed_1_0_1122_inst_req_0;
      W_condx_xend_ifx_xend238_taken_997_delayed_1_0_1122_inst_ack_0<= wack(0);
      rreq(0) <= W_condx_xend_ifx_xend238_taken_997_delayed_1_0_1122_inst_req_1;
      W_condx_xend_ifx_xend238_taken_997_delayed_1_0_1122_inst_ack_1<= rack(0);
      W_condx_xend_ifx_xend238_taken_997_delayed_1_0_1122_inst : InterlockBuffer generic map ( -- 
        name => "W_condx_xend_ifx_xend238_taken_997_delayed_1_0_1122_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => condx_xend_ifx_xend238_taken_1044,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => condx_xend_ifx_xend238_taken_997_delayed_1_0_1124,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_iNsTr_28_1010_delayed_2_0_1140_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_iNsTr_28_1010_delayed_2_0_1140_inst_req_0;
      W_iNsTr_28_1010_delayed_2_0_1140_inst_ack_0<= wack(0);
      rreq(0) <= W_iNsTr_28_1010_delayed_2_0_1140_inst_req_1;
      W_iNsTr_28_1010_delayed_2_0_1140_inst_ack_1<= rack(0);
      W_iNsTr_28_1010_delayed_2_0_1140_inst : InterlockBuffer generic map ( -- 
        name => "W_iNsTr_28_1010_delayed_2_0_1140_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_28_600,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_28_1010_delayed_2_0_1142,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_ifx_xend186_exec_guard_658_inst
    process(whilex_xbody_ifx_xend186_taken_657) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := whilex_xbody_ifx_xend186_taken_657(0 downto 0);
      ifx_xend186_exec_guard_660 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xend186_ifx_xend238_taken_668_inst
    process(ifx_xend186_exec_guard_660) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xend186_exec_guard_660(0 downto 0);
      ifx_xend186_ifx_xend238_taken_670 <= tmp_var; -- 
    end process;
    W_ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1045_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1045_inst_req_0;
      W_ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1045_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1045_inst_req_1;
      W_ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1045_inst_ack_1<= rack(0);
      W_ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1045_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1045_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend186_ifx_xend238_taken_670,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1047,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_ifx_xend253_whilex_xend_taken_1326_inst
    process(cmp284_1325) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp284_1325(0 downto 0);
      ifx_xend253_whilex_xend_taken_1328 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xend_exec_guard_671_inst
    process(whilex_xbody_ifx_xend_taken_653) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := whilex_xbody_ifx_xend_taken_653(0 downto 0);
      ifx_xend_exec_guard_673 <= tmp_var; -- 
    end process;
    W_ifx_xend_exec_guard_686_delayed_1_0_686_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend_exec_guard_686_delayed_1_0_686_inst_req_0;
      W_ifx_xend_exec_guard_686_delayed_1_0_686_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend_exec_guard_686_delayed_1_0_686_inst_req_1;
      W_ifx_xend_exec_guard_686_delayed_1_0_686_inst_ack_1<= rack(0);
      W_ifx_xend_exec_guard_686_delayed_1_0_686_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend_exec_guard_686_delayed_1_0_686_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend_exec_guard_673,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend_exec_guard_686_delayed_1_0_688,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend_exec_guard_693_delayed_1_0_696_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend_exec_guard_693_delayed_1_0_696_inst_req_0;
      W_ifx_xend_exec_guard_693_delayed_1_0_696_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend_exec_guard_693_delayed_1_0_696_inst_req_1;
      W_ifx_xend_exec_guard_693_delayed_1_0_696_inst_ack_1<= rack(0);
      W_ifx_xend_exec_guard_693_delayed_1_0_696_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend_exec_guard_693_delayed_1_0_696_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend_exec_guard_673,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend_exec_guard_693_delayed_1_0_698,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend_exec_guard_700_delayed_1_0_706_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend_exec_guard_700_delayed_1_0_706_inst_req_0;
      W_ifx_xend_exec_guard_700_delayed_1_0_706_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend_exec_guard_700_delayed_1_0_706_inst_req_1;
      W_ifx_xend_exec_guard_700_delayed_1_0_706_inst_ack_1<= rack(0);
      W_ifx_xend_exec_guard_700_delayed_1_0_706_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend_exec_guard_700_delayed_1_0_706_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend_exec_guard_673,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend_exec_guard_700_delayed_1_0_708,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend_exec_guard_705_delayed_2_0_714_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend_exec_guard_705_delayed_2_0_714_inst_req_0;
      W_ifx_xend_exec_guard_705_delayed_2_0_714_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend_exec_guard_705_delayed_2_0_714_inst_req_1;
      W_ifx_xend_exec_guard_705_delayed_2_0_714_inst_ack_1<= rack(0);
      W_ifx_xend_exec_guard_705_delayed_2_0_714_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend_exec_guard_705_delayed_2_0_714_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend_exec_guard_673,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend_exec_guard_705_delayed_2_0_716,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend_exec_guard_718_delayed_2_0_733_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend_exec_guard_718_delayed_2_0_733_inst_req_0;
      W_ifx_xend_exec_guard_718_delayed_2_0_733_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend_exec_guard_718_delayed_2_0_733_inst_req_1;
      W_ifx_xend_exec_guard_718_delayed_2_0_733_inst_ack_1<= rack(0);
      W_ifx_xend_exec_guard_718_delayed_2_0_733_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend_exec_guard_718_delayed_2_0_733_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend_exec_guard_673,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend_exec_guard_718_delayed_2_0_735,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend_exec_guard_725_delayed_2_0_743_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend_exec_guard_725_delayed_2_0_743_inst_req_0;
      W_ifx_xend_exec_guard_725_delayed_2_0_743_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend_exec_guard_725_delayed_2_0_743_inst_req_1;
      W_ifx_xend_exec_guard_725_delayed_2_0_743_inst_ack_1<= rack(0);
      W_ifx_xend_exec_guard_725_delayed_2_0_743_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend_exec_guard_725_delayed_2_0_743_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend_exec_guard_673,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend_exec_guard_725_delayed_2_0_745,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen180_exec_guard_768_delayed_6_0_792_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen180_exec_guard_768_delayed_6_0_792_inst_req_0;
      W_ifx_xthen180_exec_guard_768_delayed_6_0_792_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen180_exec_guard_768_delayed_6_0_792_inst_req_1;
      W_ifx_xthen180_exec_guard_768_delayed_6_0_792_inst_ack_1<= rack(0);
      W_ifx_xthen180_exec_guard_768_delayed_6_0_792_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen180_exec_guard_768_delayed_6_0_792_inst",
        buffer_size => 6,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen180_exec_guard_775,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen180_exec_guard_768_delayed_6_0_794,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_ifx_xthen180_exec_guard_773_inst
    process(ifx_xend_ifx_xthen180_taken_766) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xend_ifx_xthen180_taken_766(0 downto 0);
      ifx_xthen180_exec_guard_775 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xthen180_ifx_xthen191_taken_800_inst
    process(ifx_xthen180_exec_guard_775) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xthen180_exec_guard_775(0 downto 0);
      ifx_xthen180_ifx_xthen191_taken_802 <= tmp_var; -- 
    end process;
    W_ifx_xthen180_ifx_xthen191_taken_807_delayed_12_0_833_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen180_ifx_xthen191_taken_807_delayed_12_0_833_inst_req_0;
      W_ifx_xthen180_ifx_xthen191_taken_807_delayed_12_0_833_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen180_ifx_xthen191_taken_807_delayed_12_0_833_inst_req_1;
      W_ifx_xthen180_ifx_xthen191_taken_807_delayed_12_0_833_inst_ack_1<= rack(0);
      W_ifx_xthen180_ifx_xthen191_taken_807_delayed_12_0_833_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen180_ifx_xthen191_taken_807_delayed_12_0_833_inst",
        buffer_size => 12,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen180_ifx_xthen191_taken_802,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen180_ifx_xthen191_taken_807_delayed_12_0_835,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen191_condx_xend_taken_911_delayed_1_0_991_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen191_condx_xend_taken_911_delayed_1_0_991_inst_req_0;
      W_ifx_xthen191_condx_xend_taken_911_delayed_1_0_991_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen191_condx_xend_taken_911_delayed_1_0_991_inst_req_1;
      W_ifx_xthen191_condx_xend_taken_911_delayed_1_0_991_inst_ack_1<= rack(0);
      W_ifx_xthen191_condx_xend_taken_911_delayed_1_0_991_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen191_condx_xend_taken_911_delayed_1_0_991_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen191_condx_xend_taken_896,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen191_condx_xend_taken_911_delayed_1_0_993,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen191_condx_xend_taken_918_delayed_2_0_1001_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen191_condx_xend_taken_918_delayed_2_0_1001_inst_req_0;
      W_ifx_xthen191_condx_xend_taken_918_delayed_2_0_1001_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen191_condx_xend_taken_918_delayed_2_0_1001_inst_req_1;
      W_ifx_xthen191_condx_xend_taken_918_delayed_2_0_1001_inst_ack_1<= rack(0);
      W_ifx_xthen191_condx_xend_taken_918_delayed_2_0_1001_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen191_condx_xend_taken_918_delayed_2_0_1001_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen191_condx_xend_taken_896,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen191_condx_xend_taken_918_delayed_2_0_1003,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen191_exec_guard_823_delayed_1_0_856_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen191_exec_guard_823_delayed_1_0_856_inst_req_0;
      W_ifx_xthen191_exec_guard_823_delayed_1_0_856_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen191_exec_guard_823_delayed_1_0_856_inst_req_1;
      W_ifx_xthen191_exec_guard_823_delayed_1_0_856_inst_ack_1<= rack(0);
      W_ifx_xthen191_exec_guard_823_delayed_1_0_856_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen191_exec_guard_823_delayed_1_0_856_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen191_exec_guard_807,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen191_exec_guard_823_delayed_1_0_858,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen191_exec_guard_829_delayed_1_0_865_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen191_exec_guard_829_delayed_1_0_865_inst_req_0;
      W_ifx_xthen191_exec_guard_829_delayed_1_0_865_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen191_exec_guard_829_delayed_1_0_865_inst_req_1;
      W_ifx_xthen191_exec_guard_829_delayed_1_0_865_inst_ack_1<= rack(0);
      W_ifx_xthen191_exec_guard_829_delayed_1_0_865_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen191_exec_guard_829_delayed_1_0_865_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen191_exec_guard_807,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen191_exec_guard_829_delayed_1_0_867,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen191_exec_guard_838_delayed_1_0_880_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen191_exec_guard_838_delayed_1_0_880_inst_req_0;
      W_ifx_xthen191_exec_guard_838_delayed_1_0_880_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen191_exec_guard_838_delayed_1_0_880_inst_req_1;
      W_ifx_xthen191_exec_guard_838_delayed_1_0_880_inst_ack_1<= rack(0);
      W_ifx_xthen191_exec_guard_838_delayed_1_0_880_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen191_exec_guard_838_delayed_1_0_880_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen191_exec_guard_807,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen191_exec_guard_838_delayed_1_0_882,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen191_exec_guard_845_delayed_1_0_889_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen191_exec_guard_845_delayed_1_0_889_inst_req_0;
      W_ifx_xthen191_exec_guard_845_delayed_1_0_889_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen191_exec_guard_845_delayed_1_0_889_inst_req_1;
      W_ifx_xthen191_exec_guard_845_delayed_1_0_889_inst_ack_1<= rack(0);
      W_ifx_xthen191_exec_guard_845_delayed_1_0_889_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen191_exec_guard_845_delayed_1_0_889_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen191_exec_guard_807,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen191_exec_guard_845_delayed_1_0_891,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen191_exec_guard_850_delayed_1_0_897_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen191_exec_guard_850_delayed_1_0_897_inst_req_0;
      W_ifx_xthen191_exec_guard_850_delayed_1_0_897_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen191_exec_guard_850_delayed_1_0_897_inst_req_1;
      W_ifx_xthen191_exec_guard_850_delayed_1_0_897_inst_ack_1<= rack(0);
      W_ifx_xthen191_exec_guard_850_delayed_1_0_897_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen191_exec_guard_850_delayed_1_0_897_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen191_exec_guard_807,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen191_exec_guard_850_delayed_1_0_899,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_ifx_xthen247_exec_guard_1178_inst
    process(ifx_xend238_ifx_xthen247_taken_1171) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xend238_ifx_xthen247_taken_1171(0 downto 0);
      ifx_xthen247_exec_guard_1180 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xthen247_ifx_xend253_taken_1205_inst
    process(ifx_xthen247_exec_guard_1180) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xthen247_exec_guard_1180(0 downto 0);
      ifx_xthen247_ifx_xend253_taken_1207 <= tmp_var; -- 
    end process;
    W_inc265_1139_delayed_1_0_1287_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_inc265_1139_delayed_1_0_1287_inst_req_0;
      W_inc265_1139_delayed_1_0_1287_inst_ack_0<= wack(0);
      rreq(0) <= W_inc265_1139_delayed_1_0_1287_inst_req_1;
      W_inc265_1139_delayed_1_0_1287_inst_ack_1<= rack(0);
      W_inc265_1139_delayed_1_0_1287_inst : InterlockBuffer generic map ( -- 
        name => "W_inc265_1139_delayed_1_0_1287_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc265_1268,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc265_1139_delayed_1_0_1289,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_input_wordx_x1_707_delayed_2_0_717_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_input_wordx_x1_707_delayed_2_0_717_inst_req_0;
      W_input_wordx_x1_707_delayed_2_0_717_inst_ack_0<= wack(0);
      rreq(0) <= W_input_wordx_x1_707_delayed_2_0_717_inst_req_1;
      W_input_wordx_x1_707_delayed_2_0_717_inst_ack_1<= rack(0);
      W_input_wordx_x1_707_delayed_2_0_717_inst : InterlockBuffer generic map ( -- 
        name => "W_input_wordx_x1_707_delayed_2_0_717_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_wordx_x1_640,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => input_wordx_x1_707_delayed_2_0_719,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_landx_xlhsx_xtrue208_condx_xend_taken_921_delayed_1_0_1008_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue208_condx_xend_taken_921_delayed_1_0_1008_inst_req_0;
      W_landx_xlhsx_xtrue208_condx_xend_taken_921_delayed_1_0_1008_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue208_condx_xend_taken_921_delayed_1_0_1008_inst_req_1;
      W_landx_xlhsx_xtrue208_condx_xend_taken_921_delayed_1_0_1008_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue208_condx_xend_taken_921_delayed_1_0_1008_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue208_condx_xend_taken_921_delayed_1_0_1008_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue208_condx_xend_taken_942,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue208_condx_xend_taken_921_delayed_1_0_1010,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_landx_xlhsx_xtrue208_exec_guard_863_delayed_1_0_917_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue208_exec_guard_863_delayed_1_0_917_inst_req_0;
      W_landx_xlhsx_xtrue208_exec_guard_863_delayed_1_0_917_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue208_exec_guard_863_delayed_1_0_917_inst_req_1;
      W_landx_xlhsx_xtrue208_exec_guard_863_delayed_1_0_917_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue208_exec_guard_863_delayed_1_0_917_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue208_exec_guard_863_delayed_1_0_917_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue208_exec_guard_908,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue208_exec_guard_863_delayed_1_0_919,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_926_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_926_inst_req_0;
      W_landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_926_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_926_inst_req_1;
      W_landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_926_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_926_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_926_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue208_exec_guard_908,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_928,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_934_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_934_inst_req_0;
      W_landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_934_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_934_inst_req_1;
      W_landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_934_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_934_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_934_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue208_exec_guard_908,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_936,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_landx_xlhsx_xtrue208_exec_guard_906_inst
    process(ifx_xthen191_landx_xlhsx_xtrue208_taken_905) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xthen191_landx_xlhsx_xtrue208_taken_905(0 downto 0);
      landx_xlhsx_xtrue208_exec_guard_908 <= tmp_var; -- 
    end process;
    W_landx_xlhsx_xtrue219_condx_xend_taken_924_delayed_1_0_1015_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue219_condx_xend_taken_924_delayed_1_0_1015_inst_req_0;
      W_landx_xlhsx_xtrue219_condx_xend_taken_924_delayed_1_0_1015_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue219_condx_xend_taken_924_delayed_1_0_1015_inst_req_1;
      W_landx_xlhsx_xtrue219_condx_xend_taken_924_delayed_1_0_1015_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue219_condx_xend_taken_924_delayed_1_0_1015_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue219_condx_xend_taken_924_delayed_1_0_1015_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue219_condx_xend_taken_990,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue219_condx_xend_taken_924_delayed_1_0_1017,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_landx_xlhsx_xtrue219_condx_xend_taken_988_inst
    process(landx_xlhsx_xtrue219_exec_guard_945) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := landx_xlhsx_xtrue219_exec_guard_945(0 downto 0);
      landx_xlhsx_xtrue219_condx_xend_taken_990 <= tmp_var; -- 
    end process;
    W_landx_xlhsx_xtrue219_exec_guard_894_delayed_1_0_963_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue219_exec_guard_894_delayed_1_0_963_inst_req_0;
      W_landx_xlhsx_xtrue219_exec_guard_894_delayed_1_0_963_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue219_exec_guard_894_delayed_1_0_963_inst_req_1;
      W_landx_xlhsx_xtrue219_exec_guard_894_delayed_1_0_963_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue219_exec_guard_894_delayed_1_0_963_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue219_exec_guard_894_delayed_1_0_963_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue219_exec_guard_945,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue219_exec_guard_894_delayed_1_0_965,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_landx_xlhsx_xtrue219_exec_guard_900_delayed_1_0_972_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_landx_xlhsx_xtrue219_exec_guard_900_delayed_1_0_972_inst_req_0;
      W_landx_xlhsx_xtrue219_exec_guard_900_delayed_1_0_972_inst_ack_0<= wack(0);
      rreq(0) <= W_landx_xlhsx_xtrue219_exec_guard_900_delayed_1_0_972_inst_req_1;
      W_landx_xlhsx_xtrue219_exec_guard_900_delayed_1_0_972_inst_ack_1<= rack(0);
      W_landx_xlhsx_xtrue219_exec_guard_900_delayed_1_0_972_inst : InterlockBuffer generic map ( -- 
        name => "W_landx_xlhsx_xtrue219_exec_guard_900_delayed_1_0_972_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => landx_xlhsx_xtrue219_exec_guard_945,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => landx_xlhsx_xtrue219_exec_guard_900_delayed_1_0_974,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_landx_xlhsx_xtrue219_exec_guard_943_inst
    process(landx_xlhsx_xtrue208_landx_xlhsx_xtrue219_taken_933) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := landx_xlhsx_xtrue208_landx_xlhsx_xtrue219_taken_933(0 downto 0);
      landx_xlhsx_xtrue219_exec_guard_945 <= tmp_var; -- 
    end process;
    W_o0x_x1_1155_delayed_3_0_1306_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_o0x_x1_1155_delayed_3_0_1306_inst_req_0;
      W_o0x_x1_1155_delayed_3_0_1306_inst_ack_0<= wack(0);
      rreq(0) <= W_o0x_x1_1155_delayed_3_0_1306_inst_req_1;
      W_o0x_x1_1155_delayed_3_0_1306_inst_ack_1<= rack(0);
      W_o0x_x1_1155_delayed_3_0_1306_inst : InterlockBuffer generic map ( -- 
        name => "W_o0x_x1_1155_delayed_3_0_1306_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => o0x_x1_620,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => o0x_x1_1155_delayed_3_0_1308,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_o1x_x1_1134_delayed_2_0_1279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_o1x_x1_1134_delayed_2_0_1279_inst_req_0;
      W_o1x_x1_1134_delayed_2_0_1279_inst_ack_0<= wack(0);
      rreq(0) <= W_o1x_x1_1134_delayed_2_0_1279_inst_req_1;
      W_o1x_x1_1134_delayed_2_0_1279_inst_ack_1<= rack(0);
      W_o1x_x1_1134_delayed_2_0_1279_inst : InterlockBuffer generic map ( -- 
        name => "W_o1x_x1_1134_delayed_2_0_1279_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => o1x_x1_625,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => o1x_x1_1134_delayed_2_0_1281,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_o1x_x1_860_delayed_1_0_909_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_o1x_x1_860_delayed_1_0_909_inst_req_0;
      W_o1x_x1_860_delayed_1_0_909_inst_ack_0<= wack(0);
      rreq(0) <= W_o1x_x1_860_delayed_1_0_909_inst_req_1;
      W_o1x_x1_860_delayed_1_0_909_inst_ack_1<= rack(0);
      W_o1x_x1_860_delayed_1_0_909_inst : InterlockBuffer generic map ( -- 
        name => "W_o1x_x1_860_delayed_1_0_909_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => o1x_x1_625,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => o1x_x1_860_delayed_1_0_911,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_o2x_x1_885_delayed_2_0_946_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_o2x_x1_885_delayed_2_0_946_inst_req_0;
      W_o2x_x1_885_delayed_2_0_946_inst_ack_0<= wack(0);
      rreq(0) <= W_o2x_x1_885_delayed_2_0_946_inst_req_1;
      W_o2x_x1_885_delayed_2_0_946_inst_ack_1<= rack(0);
      W_o2x_x1_885_delayed_2_0_946_inst : InterlockBuffer generic map ( -- 
        name => "W_o2x_x1_885_delayed_2_0_946_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => o2x_x1_630,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => o2x_x1_885_delayed_2_0_948,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_byte_countx_x0_1017_delayed_2_0_1150_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_byte_countx_x0_1017_delayed_2_0_1150_inst_req_0;
      W_output_byte_countx_x0_1017_delayed_2_0_1150_inst_ack_0<= wack(0);
      rreq(0) <= W_output_byte_countx_x0_1017_delayed_2_0_1150_inst_req_1;
      W_output_byte_countx_x0_1017_delayed_2_0_1150_inst_ack_1<= rack(0);
      W_output_byte_countx_x0_1017_delayed_2_0_1150_inst : InterlockBuffer generic map ( -- 
        name => "W_output_byte_countx_x0_1017_delayed_2_0_1150_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_byte_countx_x0_610,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_byte_countx_x0_1017_delayed_2_0_1152,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_shl169_728_delayed_2_0_746_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_shl169_728_delayed_2_0_746_inst_req_0;
      W_shl169_728_delayed_2_0_746_inst_ack_0<= wack(0);
      rreq(0) <= W_shl169_728_delayed_2_0_746_inst_req_1;
      W_shl169_728_delayed_2_0_746_inst_ack_1<= rack(0);
      W_shl169_728_delayed_2_0_746_inst : InterlockBuffer generic map ( -- 
        name => "W_shl169_728_delayed_2_0_746_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl169_732,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => shl169_728_delayed_2_0_748,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_target_out_offsetx_x1_890_delayed_2_0_954_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_target_out_offsetx_x1_890_delayed_2_0_954_inst_req_0;
      W_target_out_offsetx_x1_890_delayed_2_0_954_inst_ack_0<= wack(0);
      rreq(0) <= W_target_out_offsetx_x1_890_delayed_2_0_954_inst_req_1;
      W_target_out_offsetx_x1_890_delayed_2_0_954_inst_ack_1<= rack(0);
      W_target_out_offsetx_x1_890_delayed_2_0_954_inst : InterlockBuffer generic map ( -- 
        name => "W_target_out_offsetx_x1_890_delayed_2_0_954_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => target_out_offsetx_x1_595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => target_out_offsetx_x1_890_delayed_2_0_956,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_target_out_offsetx_x1_904_delayed_3_0_978_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_target_out_offsetx_x1_904_delayed_3_0_978_inst_req_0;
      W_target_out_offsetx_x1_904_delayed_3_0_978_inst_ack_0<= wack(0);
      rreq(0) <= W_target_out_offsetx_x1_904_delayed_3_0_978_inst_req_1;
      W_target_out_offsetx_x1_904_delayed_3_0_978_inst_ack_1<= rack(0);
      W_target_out_offsetx_x1_904_delayed_3_0_978_inst : InterlockBuffer generic map ( -- 
        name => "W_target_out_offsetx_x1_904_delayed_3_0_978_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => target_out_offsetx_x1_595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => target_out_offsetx_x1_904_delayed_3_0_980,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_whilex_xbody_ifx_xend_taken_651_inst
    process(cmp158_650) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp158_650(0 downto 0);
      whilex_xbody_ifx_xend_taken_653 <= tmp_var; -- 
    end process;
    addr_of_1188_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1188_final_reg_req_0;
      addr_of_1188_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1188_final_reg_req_1;
      addr_of_1188_final_reg_ack_1<= rack(0);
      addr_of_1188_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1188_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 15,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1187_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx250_1189,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1522_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1522_final_reg_req_0;
      addr_of_1522_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1522_final_reg_req_1;
      addr_of_1522_final_reg_ack_1<= rack(0);
      addr_of_1522_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1522_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 15,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1521_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx375_1523,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_284_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_284_final_reg_req_0;
      addr_of_284_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_284_final_reg_req_1;
      addr_of_284_final_reg_ack_1<= rack(0);
      addr_of_284_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_284_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 15,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_283_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_285,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_790_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_790_final_reg_req_0;
      addr_of_790_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_790_final_reg_req_1;
      addr_of_790_final_reg_ack_1<= rack(0);
      addr_of_790_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_790_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 15,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_789_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx184_791,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    input_wordx_x1_at_entry_583_644_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= input_wordx_x1_at_entry_583_644_buf_req_0;
      input_wordx_x1_at_entry_583_644_buf_ack_0<= wack(0);
      rreq(0) <= input_wordx_x1_at_entry_583_644_buf_req_1;
      input_wordx_x1_at_entry_583_644_buf_ack_1<= rack(0);
      input_wordx_x1_at_entry_583_644_buf : InterlockBuffer generic map ( -- 
        name => "input_wordx_x1_at_entry_583_644_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_wordx_x1_at_entry_583,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => input_wordx_x1_at_entry_583_644_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    target_out_offsetx_x1_at_entry_539_599_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= target_out_offsetx_x1_at_entry_539_599_buf_req_0;
      target_out_offsetx_x1_at_entry_539_599_buf_ack_0<= wack(0);
      rreq(0) <= target_out_offsetx_x1_at_entry_539_599_buf_req_1;
      target_out_offsetx_x1_at_entry_539_599_buf_ack_1<= rack(0);
      target_out_offsetx_x1_at_entry_539_599_buf : InterlockBuffer generic map ( -- 
        name => "target_out_offsetx_x1_at_entry_539_599_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => target_out_offsetx_x1_at_entry_539,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => target_out_offsetx_x1_at_entry_539_599_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1006_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1006_inst_req_0;
      type_cast_1006_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1006_inst_req_1;
      type_cast_1006_inst_ack_1<= rack(0);
      type_cast_1006_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1006_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => target_out_offsetx_x1_595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_920_920_delayed_3_0_1007,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_100_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_100_inst_req_0;
      type_cast_100_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_100_inst_req_1;
      type_cast_100_inst_ack_1<= rack(0);
      type_cast_100_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_100_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_97,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_101,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1013_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1013_inst_req_0;
      type_cast_1013_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1013_inst_req_1;
      type_cast_1013_inst_ack_1<= rack(0);
      type_cast_1013_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1013_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => target_out_offsetx_x1_595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_923_923_delayed_3_0_1014,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1025_inst
    process(add234x_xtarget_out_offsetx_x1_987) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add234x_xtarget_out_offsetx_x1_987(31 downto 0);
      type_cast_1025_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1059_inst
    process(input_wordx_x1_640) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := input_wordx_x1_640(63 downto 0);
      type_cast_1059_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1067_inst
    process(input_wordx_x0x_xph_850) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := input_wordx_x0x_xph_850(63 downto 0);
      type_cast_1067_wire <= tmp_var; -- 
    end process;
    type_cast_1073_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1073_inst_req_0;
      type_cast_1073_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1073_inst_req_1;
      type_cast_1073_inst_ack_1<= rack(0);
      type_cast_1073_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1073_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_byte_countx_x2x_xph_832,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_963_963_delayed_2_0_1074,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1078_inst
    process(input_byte_countx_x1_615) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := input_byte_countx_x1_615(7 downto 0);
      type_cast_1078_wire <= tmp_var; -- 
    end process;
    type_cast_1091_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1091_inst_req_0;
      type_cast_1091_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1091_inst_req_1;
      type_cast_1091_inst_ack_1<= rack(0);
      type_cast_1091_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1091_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_srcx_x0x_xph_819,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_975_975_delayed_2_0_1092,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1096_inst
    process(add_srcx_x1_590) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_srcx_x1_590(31 downto 0);
      type_cast_1096_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1110_inst
    process(shl175_667) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := shl175_667(63 downto 0);
      type_cast_1110_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1118_inst
    process(add173_754) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := add173_754(63 downto 0);
      type_cast_1118_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1128_inst
    process(target_out_offsetx_x1_595) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := target_out_offsetx_x1_595(31 downto 0);
      type_cast_1128_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1136_inst
    process(cond_1041) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := cond_1041(31 downto 0);
      type_cast_1136_wire <= tmp_var; -- 
    end process;
    type_cast_113_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_113_inst_req_0;
      type_cast_113_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_113_inst_req_1;
      type_cast_113_inst_ack_1<= rack(0);
      type_cast_113_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_113_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_110,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_114,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1210_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1210_inst_req_0;
      type_cast_1210_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1210_inst_req_1;
      type_cast_1210_inst_ack_1<= rack(0);
      type_cast_1210_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1210_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x1_605,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1073_1073_delayed_2_0_1211,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1215_inst
    process(inc252_1204) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := inc252_1204(31 downto 0);
      type_cast_1215_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1230_inst
    process(inc242_1159) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := inc242_1159(7 downto 0);
      type_cast_1230_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1243_inst
    process(valuex_x0448450_1121) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := valuex_x0448450_1121(63 downto 0);
      type_cast_1243_wire <= tmp_var; -- 
    end process;
    type_cast_1251_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1251_inst_req_0;
      type_cast_1251_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1251_inst_req_1;
      type_cast_1251_inst_ack_1<= rack(0);
      type_cast_1251_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1251_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => o2x_x1_630,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv257_1252,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1255_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1255_inst_req_0;
      type_cast_1255_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1255_inst_req_1;
      type_cast_1255_inst_ack_1<= rack(0);
      type_cast_1255_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1255_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub224_520,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1113_1113_delayed_2_0_1256,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1259_inst
    process(conv257_1252) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv257_1252(31 downto 0);
      type_cast_1259_wire <= tmp_var; -- 
    end process;
    type_cast_126_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_126_inst_req_0;
      type_cast_126_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_126_inst_req_1;
      type_cast_126_inst_ack_1<= rack(0);
      type_cast_126_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_126_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_122,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_127,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1271_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1271_inst_req_0;
      type_cast_1271_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1271_inst_req_1;
      type_cast_1271_inst_ack_1<= rack(0);
      type_cast_1271_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1271_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp261_1262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_41_1272,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1304_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1304_inst_req_0;
      type_cast_1304_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1304_inst_req_1;
      type_cast_1304_inst_ack_1<= rack(0);
      type_cast_1304_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1304_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp274_1301,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc278_1305,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1341_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1341_inst_req_0;
      type_cast_1341_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1341_inst_req_1;
      type_cast_1341_inst_ack_1<= rack(0);
      type_cast_1341_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1341_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1340_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv121_1342,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1349_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1349_inst_req_0;
      type_cast_1349_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1349_inst_req_1;
      type_cast_1349_inst_ack_1<= rack(0);
      type_cast_1349_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1349_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1348_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv297_1350,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1358_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1358_inst_req_0;
      type_cast_1358_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1358_inst_req_1;
      type_cast_1358_inst_ack_1<= rack(0);
      type_cast_1358_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1358_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub301_1355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv305_1359,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1368_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1368_inst_req_0;
      type_cast_1368_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1368_inst_req_1;
      type_cast_1368_inst_ack_1<= rack(0);
      type_cast_1368_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1368_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr308_1365,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv311_1369,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1378_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1378_inst_req_0;
      type_cast_1378_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1378_inst_req_1;
      type_cast_1378_inst_ack_1<= rack(0);
      type_cast_1378_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1378_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr314_1375,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv317_1379,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1388_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1388_inst_req_0;
      type_cast_1388_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1388_inst_req_1;
      type_cast_1388_inst_ack_1<= rack(0);
      type_cast_1388_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1388_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr320_1385,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv323_1389,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1398_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1398_inst_req_0;
      type_cast_1398_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1398_inst_req_1;
      type_cast_1398_inst_ack_1<= rack(0);
      type_cast_1398_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1398_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr326_1395,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv329_1399,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_139_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_139_inst_req_0;
      type_cast_139_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_139_inst_req_1;
      type_cast_139_inst_ack_1<= rack(0);
      type_cast_139_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_139_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_136,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_140,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1408_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1408_inst_req_0;
      type_cast_1408_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1408_inst_req_1;
      type_cast_1408_inst_ack_1<= rack(0);
      type_cast_1408_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1408_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr332_1405,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv335_1409,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1418_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1418_inst_req_0;
      type_cast_1418_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1418_inst_req_1;
      type_cast_1418_inst_ack_1<= rack(0);
      type_cast_1418_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1418_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr338_1415,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv341_1419,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1428_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1428_inst_req_0;
      type_cast_1428_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1428_inst_req_1;
      type_cast_1428_inst_ack_1<= rack(0);
      type_cast_1428_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1428_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr344_1425,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv347_1429,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1470_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1470_inst_req_0;
      type_cast_1470_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1470_inst_req_1;
      type_cast_1470_inst_ack_1<= rack(0);
      type_cast_1470_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1470_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_170,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp_1471,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1479_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1479_inst_req_0;
      type_cast_1479_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1479_inst_req_1;
      type_cast_1479_inst_ack_1<= rack(0);
      type_cast_1479_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1479_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_145,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp2_1480,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1513_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1513_inst_req_0;
      type_cast_1513_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1513_inst_req_1;
      type_cast_1513_inst_ack_1<= rack(0);
      type_cast_1513_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1513_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc442_1631,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1513_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_151_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_151_inst_req_0;
      type_cast_151_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_151_inst_req_1;
      type_cast_151_inst_ack_1<= rack(0);
      type_cast_151_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_151_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_148,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_152,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1530_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1530_inst_req_0;
      type_cast_1530_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1530_inst_req_1;
      type_cast_1530_inst_ack_1<= rack(0);
      type_cast_1530_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1530_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp376_1527,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv380_1531,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1540_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1540_inst_req_0;
      type_cast_1540_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1540_inst_req_1;
      type_cast_1540_inst_ack_1<= rack(0);
      type_cast_1540_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1540_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr383_1537,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv386_1541,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1550_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1550_inst_req_0;
      type_cast_1550_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1550_inst_req_1;
      type_cast_1550_inst_ack_1<= rack(0);
      type_cast_1550_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1550_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr389_1547,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv392_1551,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1560_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1560_inst_req_0;
      type_cast_1560_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1560_inst_req_1;
      type_cast_1560_inst_ack_1<= rack(0);
      type_cast_1560_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1560_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr395_1557,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv398_1561,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1570_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1570_inst_req_0;
      type_cast_1570_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1570_inst_req_1;
      type_cast_1570_inst_ack_1<= rack(0);
      type_cast_1570_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1570_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr401_1567,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv404_1571,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1580_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1580_inst_req_0;
      type_cast_1580_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1580_inst_req_1;
      type_cast_1580_inst_ack_1<= rack(0);
      type_cast_1580_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1580_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr407_1577,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv410_1581,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1590_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1590_inst_req_0;
      type_cast_1590_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1590_inst_req_1;
      type_cast_1590_inst_ack_1<= rack(0);
      type_cast_1590_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1590_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr413_1587,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv416_1591,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1600_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1600_inst_req_0;
      type_cast_1600_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1600_inst_req_1;
      type_cast_1600_inst_ack_1<= rack(0);
      type_cast_1600_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1600_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr419_1597,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv422_1601,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_164_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_164_inst_req_0;
      type_cast_164_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_164_inst_req_1;
      type_cast_164_inst_ack_1<= rack(0);
      type_cast_164_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_164_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_161,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_165,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_176_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_176_inst_req_0;
      type_cast_176_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_176_inst_req_1;
      type_cast_176_inst_ack_1<= rack(0);
      type_cast_176_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_176_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_173,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_177,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_189_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_189_inst_req_0;
      type_cast_189_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_189_inst_req_1;
      type_cast_189_inst_ack_1<= rack(0);
      type_cast_189_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_189_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_186,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_190,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_208_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_208_inst_req_0;
      type_cast_208_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_208_inst_req_1;
      type_cast_208_inst_ack_1<= rack(0);
      type_cast_208_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_208_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add30_145,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_209,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_212_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_212_inst_req_0;
      type_cast_212_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_212_inst_req_1;
      type_cast_212_inst_ack_1<= rack(0);
      type_cast_212_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_212_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add39_170,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_213,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_275_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_275_inst_req_0;
      type_cast_275_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_275_inst_req_1;
      type_cast_275_inst_ack_1<= rack(0);
      type_cast_275_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_275_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_428,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_275_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_291_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_291_inst_req_0;
      type_cast_291_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_291_inst_req_1;
      type_cast_291_inst_ack_1<= rack(0);
      type_cast_291_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_291_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call72_288,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_292,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_304_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_304_inst_req_0;
      type_cast_304_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_304_inst_req_1;
      type_cast_304_inst_ack_1<= rack(0);
      type_cast_304_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_304_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call76_301,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv78_305,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_322_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_322_inst_req_0;
      type_cast_322_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_322_inst_req_1;
      type_cast_322_inst_ack_1<= rack(0);
      type_cast_322_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_322_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call82_319,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_323,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_340_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_340_inst_req_0;
      type_cast_340_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_340_inst_req_1;
      type_cast_340_inst_ack_1<= rack(0);
      type_cast_340_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_340_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call88_337,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_341,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_358_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_358_inst_req_0;
      type_cast_358_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_358_inst_req_1;
      type_cast_358_inst_ack_1<= rack(0);
      type_cast_358_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_358_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call94_355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv96_359,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_376_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_376_inst_req_0;
      type_cast_376_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_376_inst_req_1;
      type_cast_376_inst_ack_1<= rack(0);
      type_cast_376_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_376_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call100_373,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv102_377,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_394_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_394_inst_req_0;
      type_cast_394_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_394_inst_req_1;
      type_cast_394_inst_ack_1<= rack(0);
      type_cast_394_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_394_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_391,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv108_395,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_412_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_412_inst_req_0;
      type_cast_412_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_412_inst_req_1;
      type_cast_412_inst_ack_1<= rack(0);
      type_cast_412_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_412_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call112_409,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv114_413,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_50_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_50_inst_req_0;
      type_cast_50_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_50_inst_req_1;
      type_cast_50_inst_ack_1<= rack(0);
      type_cast_50_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_50_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_46,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_51,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_542_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_542_inst_req_0;
      type_cast_542_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_542_inst_req_1;
      type_cast_542_inst_ack_1<= rack(0);
      type_cast_542_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_542_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul145_478,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_542_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_586_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_586_inst_req_0;
      type_cast_586_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_586_inst_req_1;
      type_cast_586_inst_ack_1<= rack(0);
      type_cast_586_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_586_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp155_492,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_586_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_593_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_593_inst_req_0;
      type_cast_593_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_593_inst_req_1;
      type_cast_593_inst_ack_1<= rack(0);
      type_cast_593_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_593_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_srcx_x0452_1106,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_593_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_598_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_598_inst_req_0;
      type_cast_598_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_598_inst_req_1;
      type_cast_598_inst_ack_1<= rack(0);
      type_cast_598_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_598_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => target_out_offsetx_x0_1139,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_598_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_603_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_603_inst_req_0;
      type_cast_603_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_603_inst_req_1;
      type_cast_603_inst_ack_1<= rack(0);
      type_cast_603_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_603_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc240_1149,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_603_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_608_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_608_inst_req_0;
      type_cast_608_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_608_inst_req_1;
      type_cast_608_inst_ack_1<= rack(0);
      type_cast_608_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_608_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_outx_x0_1222,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_608_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_613_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_613_inst_req_0;
      type_cast_613_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_613_inst_req_1;
      type_cast_613_inst_ack_1<= rack(0);
      type_cast_613_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_613_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_byte_countx_x1_1235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_613_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_618_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_618_inst_req_0;
      type_cast_618_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_618_inst_req_1;
      type_cast_618_inst_ack_1<= rack(0);
      type_cast_618_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_618_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_byte_countx_x2454_1088,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_618_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_623_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_623_inst_req_0;
      type_cast_623_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_623_inst_req_1;
      type_cast_623_inst_ack_1<= rack(0);
      type_cast_623_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_623_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc278x_xo0x_x1_1313,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_623_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_628_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_628_inst_req_0;
      type_cast_628_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_628_inst_req_1;
      type_cast_628_inst_ack_1<= rack(0);
      type_cast_628_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_628_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => o1x_x2_1320,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_628_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_633_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_633_inst_req_0;
      type_cast_633_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_633_inst_req_1;
      type_cast_633_inst_ack_1<= rack(0);
      type_cast_633_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_633_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => o2x_x0_1296,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_633_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_638_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_638_inst_req_0;
      type_cast_638_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_638_inst_req_1;
      type_cast_638_inst_ack_1<= rack(0);
      type_cast_638_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_638_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => valuex_x2_1248,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_638_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_63_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_63_inst_req_0;
      type_cast_63_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_63_inst_req_1;
      type_cast_63_inst_ack_1<= rack(0);
      type_cast_63_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_63_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_60,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_64,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_643_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_643_inst_req_0;
      type_cast_643_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_643_inst_req_1;
      type_cast_643_inst_ack_1<= rack(0);
      type_cast_643_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_643_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_wordx_x0456_1070,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_643_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_684_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_684_inst_req_0;
      type_cast_684_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_684_inst_req_1;
      type_cast_684_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xend_exec_guard_673(0);
      type_cast_684_inst_gI: SplitGuardInterface generic map(name => "type_cast_684_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_684_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_684_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_byte_countx_x1_615,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv163_685,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_712_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_712_inst_req_0;
      type_cast_712_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_712_inst_req_1;
      type_cast_712_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xend_exec_guard_700_delayed_1_0_708(0);
      type_cast_712_inst_gI: SplitGuardInterface generic map(name => "type_cast_712_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_712_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_712_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub165_705,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => sh_prom_713,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_75_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_75_inst_req_0;
      type_cast_75_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_75_inst_req_1;
      type_cast_75_inst_ack_1<= rack(0);
      type_cast_75_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_75_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_72,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_76,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_811_inst
    process(add182_782) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add182_782(31 downto 0);
      type_cast_811_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_814_inst
    process(add_srcx_x1_590) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := add_srcx_x1_590(31 downto 0);
      type_cast_814_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_827_inst
    process(inc162_680) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := inc162_680(7 downto 0);
      type_cast_827_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_839_inst
    process(input_wordx_x1_640) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := input_wordx_x1_640(63 downto 0);
      type_cast_839_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_847_inst
    process(tmp185_799) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp185_799(63 downto 0);
      type_cast_847_wire <= tmp_var; -- 
    end process;
    type_cast_854_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_854_inst_req_0;
      type_cast_854_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_854_inst_req_1;
      type_cast_854_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xthen191_exec_guard_807(0);
      type_cast_854_inst_gI: SplitGuardInterface generic map(name => "type_cast_854_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_854_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_854_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => o0x_x1_620,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv193_855,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_871_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_871_inst_req_0;
      type_cast_871_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_871_inst_req_1;
      type_cast_871_inst_ack_1<= rack(0);
      type_cast_871_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_871_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub205_503,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_835_835_delayed_1_0_872,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_876_inst
    process(conv193_855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv193_855(31 downto 0);
      type_cast_876_wire <= tmp_var; -- 
    end process;
    type_cast_88_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_88_inst_req_0;
      type_cast_88_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_88_inst_req_1;
      type_cast_88_inst_ack_1<= rack(0);
      type_cast_88_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_88_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_85,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_89,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_915_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_915_inst_req_0;
      type_cast_915_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_915_inst_req_1;
      type_cast_915_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  landx_xlhsx_xtrue208_exec_guard_908(0);
      type_cast_915_inst_gI: SplitGuardInterface generic map(name => "type_cast_915_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_915_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_915_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => o1x_x1_860_delayed_1_0_911,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv210_916,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_952_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_952_inst_req_0;
      type_cast_952_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_952_inst_req_1;
      type_cast_952_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  landx_xlhsx_xtrue219_exec_guard_945(0);
      type_cast_952_inst_gI: SplitGuardInterface generic map(name => "type_cast_952_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_952_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_952_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => o2x_x1_885_delayed_2_0_948,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv221_953,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1187_index_2_rename
    process(R_add_outx_x1_1186_resized) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_add_outx_x1_1186_resized;
      ov(14 downto 0) := iv;
      R_add_outx_x1_1186_scaled <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1187_index_2_resize
    process(add_outx_x1_605) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add_outx_x1_605;
      ov := iv(14 downto 0);
      R_add_outx_x1_1186_resized <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1187_root_address_inst
    process(array_obj_ref_1187_final_offset) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1187_final_offset;
      ov(14 downto 0) := iv;
      array_obj_ref_1187_root_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1521_index_2_rename
    process(R_ix_x1460_1520_resized) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x1460_1520_resized;
      ov(14 downto 0) := iv;
      R_ix_x1460_1520_scaled <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1521_index_2_resize
    process(ix_x1460_1507) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x1460_1507;
      ov := iv(14 downto 0);
      R_ix_x1460_1520_resized <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1521_root_address_inst
    process(array_obj_ref_1521_final_offset) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1521_final_offset;
      ov(14 downto 0) := iv;
      array_obj_ref_1521_root_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_283_index_2_rename
    process(R_ix_x0463_282_resized) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0463_282_resized;
      ov(14 downto 0) := iv;
      R_ix_x0463_282_scaled <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_283_index_2_resize
    process(ix_x0463_269) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0463_269;
      ov := iv(14 downto 0);
      R_ix_x0463_282_resized <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_283_root_address_inst
    process(array_obj_ref_283_final_offset) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_283_final_offset;
      ov(14 downto 0) := iv;
      array_obj_ref_283_root_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_789_index_2_rename
    process(R_add182_788_resized) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_add182_788_resized;
      ov(14 downto 0) := iv;
      R_add182_788_scaled <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_789_index_2_resize
    process(add182_782) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add182_782;
      ov := iv(14 downto 0);
      R_add182_788_resized <= ov(14 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_789_root_address_inst
    process(array_obj_ref_789_final_offset) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_789_final_offset;
      ov(14 downto 0) := iv;
      array_obj_ref_789_root_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1192_addr_0
    process(ptr_deref_1192_root_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1192_root_address;
      ov(14 downto 0) := iv;
      ptr_deref_1192_word_address_0 <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1192_base_resize
    process(arrayidx250_1189) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx250_1189;
      ov := iv(14 downto 0);
      ptr_deref_1192_resized_base_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1192_gather_scatter
    process(valuex_x0448450_1121) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := valuex_x0448450_1121;
      ov(63 downto 0) := iv;
      ptr_deref_1192_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1192_root_address_inst
    process(ptr_deref_1192_resized_base_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1192_resized_base_address;
      ov(14 downto 0) := iv;
      ptr_deref_1192_root_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1526_addr_0
    process(ptr_deref_1526_root_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1526_root_address;
      ov(14 downto 0) := iv;
      ptr_deref_1526_word_address_0 <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1526_base_resize
    process(arrayidx375_1523) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx375_1523;
      ov := iv(14 downto 0);
      ptr_deref_1526_resized_base_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1526_gather_scatter
    process(ptr_deref_1526_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1526_data_0;
      ov(63 downto 0) := iv;
      tmp376_1527 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1526_root_address_inst
    process(ptr_deref_1526_resized_base_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1526_resized_base_address;
      ov(14 downto 0) := iv;
      ptr_deref_1526_root_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_420_addr_0
    process(ptr_deref_420_root_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_420_root_address;
      ov(14 downto 0) := iv;
      ptr_deref_420_word_address_0 <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_420_base_resize
    process(arrayidx_285) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_285;
      ov := iv(14 downto 0);
      ptr_deref_420_resized_base_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_420_gather_scatter
    process(add115_418) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add115_418;
      ov(63 downto 0) := iv;
      ptr_deref_420_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_420_root_address_inst
    process(ptr_deref_420_resized_base_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_420_resized_base_address;
      ov(14 downto 0) := iv;
      ptr_deref_420_root_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_491_addr_0
    process(ptr_deref_491_root_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_491_root_address;
      ov(14 downto 0) := iv;
      ptr_deref_491_word_address_0 <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_491_base_resize
    process(iNsTr_16_488) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_16_488;
      ov := iv(14 downto 0);
      ptr_deref_491_resized_base_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_491_gather_scatter
    process(ptr_deref_491_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_491_data_0;
      ov(63 downto 0) := iv;
      tmp155_492 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_491_root_address_inst
    process(ptr_deref_491_resized_base_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_491_resized_base_address;
      ov(14 downto 0) := iv;
      ptr_deref_491_root_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_798_addr_0
    process(ptr_deref_798_root_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_798_root_address;
      ov(14 downto 0) := iv;
      ptr_deref_798_word_address_0 <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_798_base_resize
    process(arrayidx184_791) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx184_791;
      ov := iv(14 downto 0);
      ptr_deref_798_resized_base_address <= ov(14 downto 0);
      --
    end process;
    -- equivalence ptr_deref_798_gather_scatter
    process(ptr_deref_798_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_798_data_0;
      ov(63 downto 0) := iv;
      tmp185_799 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_798_root_address_inst
    process(ptr_deref_798_resized_base_address) --
      variable iv : std_logic_vector(14 downto 0);
      variable ov : std_logic_vector(14 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_798_resized_base_address;
      ov(14 downto 0) := iv;
      ptr_deref_798_root_address <= ov(14 downto 0);
      --
    end process;
    do_while_stmt_588_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1331_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_588_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_588_branch_req_0,
          ack0 => do_while_stmt_588_branch_ack_0,
          ack1 => do_while_stmt_588_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1332_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ifx_xend253_whilex_xend_taken_1328;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1332_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1332_branch_req_0,
          ack0 => if_stmt_1332_branch_ack_0,
          ack1 => if_stmt_1332_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1461_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp369459_1460;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1461_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1461_branch_req_0,
          ack0 => if_stmt_1461_branch_ack_0,
          ack1 => if_stmt_1461_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1637_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond7_1636;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1637_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1637_branch_req_0,
          ack0 => if_stmt_1637_branch_ack_0,
          ack1 => if_stmt_1637_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_231_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp462_230;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_231_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_231_branch_req_0,
          ack0 => if_stmt_231_branch_ack_0,
          ack1 => if_stmt_231_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_434_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_433;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_434_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_434_branch_req_0,
          ack0 => if_stmt_434_branch_ack_0,
          ack1 => if_stmt_434_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1267_inst
    process(o2x_x1_630) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(o2x_x1_630, type_cast_1266_wire_constant, tmp_var);
      inc265_1268 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1285_inst
    process(inc268_1278, o1x_x1_1134_delayed_2_0_1281) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc268_1278, o1x_x1_1134_delayed_2_0_1281, tmp_var);
      o1x_x0_1286 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1312_inst
    process(inc278_1305, o0x_x1_1155_delayed_3_0_1308) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc278_1305, o0x_x1_1155_delayed_3_0_1308, tmp_var);
      inc278x_xo0x_x1_1313 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1040_inst
    process(condx_xin_1031) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(condx_xin_1031, type_cast_1039_wire_constant, tmp_var);
      cond_1041 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1148_inst
    process(iNsTr_28_1010_delayed_2_0_1142) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_28_1010_delayed_2_0_1142, type_cast_1147_wire_constant, tmp_var);
      inc240_1149 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1203_inst
    process(add_outx_x1_1059_delayed_2_0_1197) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_outx_x1_1059_delayed_2_0_1197, type_cast_1202_wire_constant, tmp_var);
      inc252_1204 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1630_inst
    process(ix_x1460_1507) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ix_x1460_1507, type_cast_1629_wire_constant, tmp_var);
      inc442_1631 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_427_inst
    process(ix_x0463_269) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ix_x0463_269, type_cast_426_wire_constant, tmp_var);
      inc_428 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_472_inst
    process(mul143_468, conv138_463) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul143_468, conv138_463, tmp_var);
      add144_473 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_497_inst
    process(conv61_209) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv61_209, type_cast_496_wire_constant, tmp_var);
      sub204_498 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_508_inst
    process(conv63_213) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv63_213, type_cast_507_wire_constant, tmp_var);
      sub215_509 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_519_inst
    process(add48_195) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add48_195, type_cast_518_wire_constant, tmp_var);
      sub224_520 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_781_inst
    process(add_srcx_x1_590) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_srcx_x1_590, type_cast_780_wire_constant, tmp_var);
      add182_782 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_961_inst
    process(target_out_offsetx_x1_890_delayed_2_0_956, mul233_531) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(target_out_offsetx_x1_890_delayed_2_0_956, mul233_531, tmp_var);
      add234_962 <= tmp_var; --
    end process;
    -- binary operator ADD_u8_u8_1158_inst
    process(output_byte_countx_x0_1017_delayed_2_0_1152) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(output_byte_countx_x0_1017_delayed_2_0_1152, type_cast_1157_wire_constant, tmp_var);
      inc242_1159 <= tmp_var; --
    end process;
    -- binary operator ADD_u8_u8_679_inst
    process(input_byte_countx_x1_615) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_byte_countx_x1_615, type_cast_678_wire_constant, tmp_var);
      inc162_680 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1170_inst
    process(ifx_xend238_exec_guard_1052, cmp245_1166) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ifx_xend238_exec_guard_1052, cmp245_1166, tmp_var);
      ifx_xend238_ifx_xthen247_taken_1171 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1176_inst
    process(ifx_xend238_exec_guard_1052, NOT_u1_u1_1175_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ifx_xend238_exec_guard_1052, NOT_u1_u1_1175_wire, tmp_var);
      ifx_xend238_ifx_xend253_taken_1177 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_765_inst
    process(ifx_xend_exec_guard_673, cmp178_761) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ifx_xend_exec_guard_673, cmp178_761, tmp_var);
      ifx_xend_ifx_xthen180_taken_766 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_771_inst
    process(ifx_xend_exec_guard_673, NOT_u1_u1_770_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ifx_xend_exec_guard_673, NOT_u1_u1_770_wire, tmp_var);
      ifx_xend_ifx_xthen191_taken_772 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_895_inst
    process(ifx_xthen191_exec_guard_845_delayed_1_0_891, orx_xcond_888) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ifx_xthen191_exec_guard_845_delayed_1_0_891, orx_xcond_888, tmp_var);
      ifx_xthen191_condx_xend_taken_896 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_904_inst
    process(ifx_xthen191_exec_guard_850_delayed_1_0_899, NOT_u1_u1_903_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ifx_xthen191_exec_guard_850_delayed_1_0_899, NOT_u1_u1_903_wire, tmp_var);
      ifx_xthen191_landx_xlhsx_xtrue208_taken_905 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_932_inst
    process(landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_928, cmp217_925) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(landx_xlhsx_xtrue208_exec_guard_870_delayed_1_0_928, cmp217_925, tmp_var);
      landx_xlhsx_xtrue208_landx_xlhsx_xtrue219_taken_933 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_941_inst
    process(landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_936, NOT_u1_u1_940_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(landx_xlhsx_xtrue208_exec_guard_875_delayed_1_0_936, NOT_u1_u1_940_wire, tmp_var);
      landx_xlhsx_xtrue208_condx_xend_taken_942 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_462_inst
    process(shr130444_457) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr130444_457, type_cast_461_wire_constant, tmp_var);
      conv138_463 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_525_inst
    process(sub_451) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(sub_451, type_cast_524_wire_constant, tmp_var);
      mul230_526 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_741_inst
    process(shr166_725) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(shr166_725, type_cast_740_wire_constant, tmp_var);
      conv172445_742 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1300_inst
    process(o1x_x0_1286, add39_170) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(o1x_x0_1286, add39_170, tmp_var);
      cmp274_1301 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1324_inst
    process(inc278x_xo0x_x1_1313, add30_145) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc278x_xo0x_x1_1313, add30_145, tmp_var);
      cmp284_1325 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1635_inst
    process(inc442_1631, umax6_1504) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc442_1631, umax6_1504, tmp_var);
      exitcond7_1636 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_432_inst
    process(inc_428, umax_266) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_428, umax_266, tmp_var);
      exitcond_433 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_649_inst
    process(iNsTr_28_600, target_out_offsetx_x1_595) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(iNsTr_28_600, target_out_offsetx_x1_595, tmp_var);
      cmp158_650 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_924_inst
    process(conv210_916, sub216_514) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv210_916, sub216_514, tmp_var);
      cmp217_925 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_970_inst
    process(conv221_953, sub224_520) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv221_953, sub224_520, tmp_var);
      cmp225_971 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_1165_inst
    process(inc242_1159) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc242_1159, type_cast_1164_wire_constant, tmp_var);
      cmp245_1166 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_760_inst
    process(inc162_680) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc162_680, type_cast_759_wire_constant, tmp_var);
      cmp178_761 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1490_inst
    process(tmp3_1485) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp3_1485, type_cast_1489_wire_constant, tmp_var);
      tmp4_1491 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_252_inst
    process(tmp9_247) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_247, type_cast_251_wire_constant, tmp_var);
      tmp10_253 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_456_inst
    process(sub_451) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_451, type_cast_455_wire_constant, tmp_var);
      shr130444_457 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1364_inst
    process(sub301_1355) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub301_1355, type_cast_1363_wire_constant, tmp_var);
      shr308_1365 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1374_inst
    process(sub301_1355) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub301_1355, type_cast_1373_wire_constant, tmp_var);
      shr314_1375 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1384_inst
    process(sub301_1355) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub301_1355, type_cast_1383_wire_constant, tmp_var);
      shr320_1385 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1394_inst
    process(sub301_1355) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub301_1355, type_cast_1393_wire_constant, tmp_var);
      shr326_1395 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1404_inst
    process(sub301_1355) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub301_1355, type_cast_1403_wire_constant, tmp_var);
      shr332_1405 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1414_inst
    process(sub301_1355) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub301_1355, type_cast_1413_wire_constant, tmp_var);
      shr338_1415 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1424_inst
    process(sub301_1355) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub301_1355, type_cast_1423_wire_constant, tmp_var);
      shr344_1425 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1536_inst
    process(tmp376_1527) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1527, type_cast_1535_wire_constant, tmp_var);
      shr383_1537 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1546_inst
    process(tmp376_1527) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1527, type_cast_1545_wire_constant, tmp_var);
      shr389_1547 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1556_inst
    process(tmp376_1527) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1527, type_cast_1555_wire_constant, tmp_var);
      shr395_1557 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1566_inst
    process(tmp376_1527) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1527, type_cast_1565_wire_constant, tmp_var);
      shr401_1567 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1576_inst
    process(tmp376_1527) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1527, type_cast_1575_wire_constant, tmp_var);
      shr407_1577 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1586_inst
    process(tmp376_1527) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1527, type_cast_1585_wire_constant, tmp_var);
      shr413_1587 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1596_inst
    process(tmp376_1527) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp376_1527, type_cast_1595_wire_constant, tmp_var);
      shr419_1597 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_724_inst
    process(input_wordx_x1_707_delayed_2_0_719, sh_prom_713) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(input_wordx_x1_707_delayed_2_0_719, sh_prom_713, tmp_var);
      shr166_725 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1475_inst
    process(add48_195, tmp_1471) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add48_195, tmp_1471, tmp_var);
      tmp1_1476 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1484_inst
    process(tmp1_1476, tmp2_1480) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_1476, tmp2_1480, tmp_var);
      tmp3_1485 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_199_inst
    process(add12_94, add_69) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add12_94, add_69, tmp_var);
      mul_200 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_204_inst
    process(mul_200, add21_119) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_200, add21_119, tmp_var);
      mul58_205 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_217_inst
    process(conv63_213, conv61_209) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv63_213, conv61_209, tmp_var);
      mul64_218 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_222_inst
    process(mul64_218, add48_195) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul64_218, add48_195, tmp_var);
      mul67_223 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_241_inst
    process(add12_94, add_69) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add12_94, add_69, tmp_var);
      tmp8_242 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_246_inst
    process(tmp8_242, add21_119) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp8_242, add21_119, tmp_var);
      tmp9_247 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_467_inst
    process(conv138_463, conv63_213) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv138_463, conv63_213, tmp_var);
      mul143_468 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_477_inst
    process(add144_473, add48_195) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add144_473, add48_195, tmp_var);
      mul145_478 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_530_inst
    process(mul230_526, add21_119) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul230_526, add21_119, tmp_var);
      mul233_531 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1175_inst
    process(cmp245_1166) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp245_1166, tmp_var);
      NOT_u1_u1_1175_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1331_inst
    process(cmp284_1325) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp284_1325, tmp_var);
      NOT_u1_u1_1331_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_656_inst
    process(cmp158_650) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp158_650, tmp_var);
      whilex_xbody_ifx_xend186_taken_657 <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_770_inst
    process(cmp178_761) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp178_761, tmp_var);
      NOT_u1_u1_770_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_903_inst
    process(orx_xcond_888) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", orx_xcond_888, tmp_var);
      NOT_u1_u1_903_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_940_inst
    process(cmp217_925) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp217_925, tmp_var);
      NOT_u1_u1_940_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u16_u16_144_inst
    process(shl27_133, conv29_140) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_133, conv29_140, tmp_var);
      add30_145 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_169_inst
    process(shl36_158, conv38_165) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_158, conv38_165, tmp_var);
      add39_170 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1051_inst
    process(condx_xend_ifx_xend238_taken_1044, ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1047) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(condx_xend_ifx_xend238_taken_1044, ifx_xend186_ifx_xend238_taken_945_delayed_2_0_1047, tmp_var);
      ifx_xend238_exec_guard_1052 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_806_inst
    process(ifx_xend_ifx_xthen191_taken_772, ifx_xthen180_ifx_xthen191_taken_802) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(ifx_xend_ifx_xthen191_taken_772, ifx_xthen180_ifx_xthen191_taken_802, tmp_var);
      ifx_xthen191_exec_guard_807 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_887_inst
    process(cmp196_864, cmp206_879) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(cmp196_864, cmp206_879, tmp_var);
      orx_xcond_888 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_998_inst
    process(landx_xlhsx_xtrue208_condx_xend_taken_942, landx_xlhsx_xtrue219_condx_xend_taken_990) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(landx_xlhsx_xtrue208_condx_xend_taken_942, landx_xlhsx_xtrue219_condx_xend_taken_990, tmp_var);
      OR_u1_u1_998_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_999_inst
    process(ifx_xthen191_condx_xend_taken_911_delayed_1_0_993, OR_u1_u1_998_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(ifx_xthen191_condx_xend_taken_911_delayed_1_0_993, OR_u1_u1_998_wire, tmp_var);
      condx_xend_exec_guard_1000 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_118_inst
    process(shl18_107, conv20_114) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_107, conv20_114, tmp_var);
      add21_119 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_194_inst
    process(shl45_183, conv47_190) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_183, conv47_190, tmp_var);
      add48_195 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_68_inst
    process(shl_57, conv3_64) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_57, conv3_64, tmp_var);
      add_69 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_93_inst
    process(shl9_82, conv11_89) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_82, conv11_89, tmp_var);
      add12_94 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_309_inst
    process(shl75_298, conv78_305) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl75_298, conv78_305, tmp_var);
      add79_310 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_327_inst
    process(shl81_316, conv84_323) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl81_316, conv84_323, tmp_var);
      add85_328 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_345_inst
    process(shl87_334, conv90_341) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl87_334, conv90_341, tmp_var);
      add91_346 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_363_inst
    process(shl93_352, conv96_359) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl93_352, conv96_359, tmp_var);
      add97_364 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_381_inst
    process(shl99_370, conv102_377) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl99_370, conv102_377, tmp_var);
      add103_382 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_399_inst
    process(shl105_388, conv108_395) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_388, conv108_395, tmp_var);
      add109_400 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_417_inst
    process(shl111_406, conv114_413) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl111_406, conv114_413, tmp_var);
      add115_418 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_753_inst
    process(conv172445_742, shl169_728_delayed_2_0_748) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv172445_742, shl169_728_delayed_2_0_748, tmp_var);
      add173_754 <= tmp_var; --
    end process;
    -- binary operator SGT_i32_u1_878_inst
    process(type_cast_876_wire, type_cast_835_835_delayed_1_0_872) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(type_cast_876_wire, type_cast_835_835_delayed_1_0_872, tmp_var);
      cmp206_879 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_132_inst
    process(conv26_127) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_127, type_cast_131_wire_constant, tmp_var);
      shl27_133 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_157_inst
    process(conv35_152) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_152, type_cast_156_wire_constant, tmp_var);
      shl36_158 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_106_inst
    process(conv17_101) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_101, type_cast_105_wire_constant, tmp_var);
      shl18_107 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_182_inst
    process(conv44_177) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_177, type_cast_181_wire_constant, tmp_var);
      shl45_183 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_56_inst
    process(conv1_51) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_51, type_cast_55_wire_constant, tmp_var);
      shl_57 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_694_inst
    process(conv163_685) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv163_685, type_cast_693_wire_constant, tmp_var);
      mul164_695 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_81_inst
    process(conv8_76) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_76, type_cast_80_wire_constant, tmp_var);
      shl9_82 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_297_inst
    process(conv73_292) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv73_292, type_cast_296_wire_constant, tmp_var);
      shl75_298 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_315_inst
    process(add79_310) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add79_310, type_cast_314_wire_constant, tmp_var);
      shl81_316 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_333_inst
    process(add85_328) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add85_328, type_cast_332_wire_constant, tmp_var);
      shl87_334 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_351_inst
    process(add91_346) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add91_346, type_cast_350_wire_constant, tmp_var);
      shl93_352 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_369_inst
    process(add97_364) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add97_364, type_cast_368_wire_constant, tmp_var);
      shl99_370 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_387_inst
    process(add103_382) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add103_382, type_cast_386_wire_constant, tmp_var);
      shl105_388 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_405_inst
    process(add109_400) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add109_400, type_cast_404_wire_constant, tmp_var);
      shl111_406 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_666_inst
    process(valuex_x1_635) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(valuex_x1_635, type_cast_665_wire_constant, tmp_var);
      shl175_667 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_731_inst
    process(valuex_x1_635) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(valuex_x1_635, type_cast_730_wire_constant, tmp_var);
      shl169_732 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1261_inst
    process(type_cast_1259_wire, type_cast_1113_1113_delayed_2_0_1256) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1259_wire, type_cast_1113_1113_delayed_2_0_1256, tmp_var);
      cmp261_1262 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_450_inst
    process(conv61_209, add_69) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv61_209, add_69, tmp_var);
      sub_451 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_502_inst
    process(sub204_498, conv138_463) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(sub204_498, conv138_463, tmp_var);
      sub205_503 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_513_inst
    process(sub215_509, conv138_463) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(sub215_509, conv138_463, tmp_var);
      sub216_514 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_704_inst
    process(type_cast_702_wire_constant, mul164_695) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(type_cast_702_wire_constant, mul164_695, tmp_var);
      sub165_705 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1354_inst
    process(conv297_1350, conv121_1342) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv297_1350, conv121_1342, tmp_var);
      sub301_1355 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1459_inst
    process(mul67_223) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul67_223, type_cast_1458_wire_constant, tmp_var);
      cmp369459_1460 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1496_inst
    process(tmp4_1491) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp4_1491, type_cast_1495_wire_constant, tmp_var);
      tmp5_1497 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_228_inst
    process(mul58_205) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul58_205, type_cast_227_wire_constant, tmp_var);
      cmp462_230 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_258_inst
    process(tmp10_253) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp10_253, type_cast_257_wire_constant, tmp_var);
      tmp11_259 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_863_inst
    process(conv193_855, conv138_463) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(conv193_855, conv138_463, tmp_var);
      cmp196_864 <= tmp_var; --
    end process;
    -- binary operator XOR_u16_u16_1277_inst
    process(iNsTr_41_1272) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntXor_proc(iNsTr_41_1272, type_cast_1276_wire_constant, tmp_var);
      inc268_1278 <= tmp_var; --
    end process;
    -- shared split operator group (119) : array_obj_ref_1187_index_offset 
    ApIntAdd_group_119: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_add_outx_x1_1186_scaled;
      array_obj_ref_1187_final_offset <= data_out(14 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1187_index_offset_req_0;
      array_obj_ref_1187_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1187_index_offset_req_1;
      array_obj_ref_1187_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_119_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_119_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_119",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 15,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 15,
          constant_operand => "100000000000000",
          constant_width => 15,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 119
    -- shared split operator group (120) : array_obj_ref_1521_index_offset 
    ApIntAdd_group_120: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x1460_1520_scaled;
      array_obj_ref_1521_final_offset <= data_out(14 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1521_index_offset_req_0;
      array_obj_ref_1521_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1521_index_offset_req_1;
      array_obj_ref_1521_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_120_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_120_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_120",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 15,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 15,
          constant_operand => "100000000000000",
          constant_width => 15,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 120
    -- shared split operator group (121) : array_obj_ref_283_index_offset 
    ApIntAdd_group_121: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0463_282_scaled;
      array_obj_ref_283_final_offset <= data_out(14 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_283_index_offset_req_0;
      array_obj_ref_283_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_283_index_offset_req_1;
      array_obj_ref_283_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_121_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_121_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_121",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 15,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 15,
          constant_operand => "000000000000000",
          constant_width => 15,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 121
    -- shared split operator group (122) : array_obj_ref_789_index_offset 
    ApIntAdd_group_122: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_add182_788_scaled;
      array_obj_ref_789_final_offset <= data_out(14 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_789_index_offset_req_0;
      array_obj_ref_789_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_789_index_offset_req_1;
      array_obj_ref_789_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_122_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_122_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_122",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 15,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 15,
          constant_operand => "000000000000000",
          constant_width => 15,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 122
    -- unary operator type_cast_1340_inst
    process(call120_445) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call120_445, tmp_var);
      type_cast_1340_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1348_inst
    process(call296_1345) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call296_1345, tmp_var);
      type_cast_1348_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_798_load_0 ptr_deref_491_load_0 ptr_deref_1526_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(44 downto 0);
      signal data_out: std_logic_vector(191 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 2, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 2, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => true);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 6);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_798_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_491_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1526_load_0_req_0;
      ptr_deref_798_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_491_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1526_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_798_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_491_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1526_load_0_req_1;
      ptr_deref_798_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_491_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1526_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <= ifx_xthen180_exec_guard_768_delayed_6_0_794(0);
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_798_word_address_0 & ptr_deref_491_word_address_0 & ptr_deref_1526_word_address_0;
      ptr_deref_798_data_0 <= data_out(191 downto 128);
      ptr_deref_491_data_0 <= data_out(127 downto 64);
      ptr_deref_1526_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 15,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(14 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1192_store_0 ptr_deref_420_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(29 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 15, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 6);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1192_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_420_store_0_req_0;
      ptr_deref_1192_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_420_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1192_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_420_store_0_req_1;
      ptr_deref_1192_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_420_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <= ifx_xthen247_exec_guard_1180(0);
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1192_word_address_0 & ptr_deref_420_word_address_0;
      data_in <= ptr_deref_1192_data_0 & ptr_deref_420_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 15,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(14 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Zeropad_input_pipe_45_inst RPIPE_Zeropad_input_pipe_135_inst RPIPE_Zeropad_input_pipe_96_inst RPIPE_Zeropad_input_pipe_59_inst RPIPE_Zeropad_input_pipe_121_inst RPIPE_Zeropad_input_pipe_109_inst RPIPE_Zeropad_input_pipe_71_inst RPIPE_Zeropad_input_pipe_84_inst RPIPE_Zeropad_input_pipe_147_inst RPIPE_Zeropad_input_pipe_160_inst RPIPE_Zeropad_input_pipe_172_inst RPIPE_Zeropad_input_pipe_185_inst RPIPE_Zeropad_input_pipe_287_inst RPIPE_Zeropad_input_pipe_300_inst RPIPE_Zeropad_input_pipe_318_inst RPIPE_Zeropad_input_pipe_336_inst RPIPE_Zeropad_input_pipe_354_inst RPIPE_Zeropad_input_pipe_372_inst RPIPE_Zeropad_input_pipe_390_inst RPIPE_Zeropad_input_pipe_408_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(159 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 19 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 19 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 19 downto 0);
      signal guard_vector : std_logic_vector( 19 downto 0);
      constant outBUFs : IntegerArray(19 downto 0) := (19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(19 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false);
      constant guardBuffering: IntegerArray(19 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2);
      -- 
    begin -- 
      reqL_unguarded(19) <= RPIPE_Zeropad_input_pipe_45_inst_req_0;
      reqL_unguarded(18) <= RPIPE_Zeropad_input_pipe_135_inst_req_0;
      reqL_unguarded(17) <= RPIPE_Zeropad_input_pipe_96_inst_req_0;
      reqL_unguarded(16) <= RPIPE_Zeropad_input_pipe_59_inst_req_0;
      reqL_unguarded(15) <= RPIPE_Zeropad_input_pipe_121_inst_req_0;
      reqL_unguarded(14) <= RPIPE_Zeropad_input_pipe_109_inst_req_0;
      reqL_unguarded(13) <= RPIPE_Zeropad_input_pipe_71_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Zeropad_input_pipe_84_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Zeropad_input_pipe_147_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Zeropad_input_pipe_160_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Zeropad_input_pipe_172_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Zeropad_input_pipe_185_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Zeropad_input_pipe_287_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Zeropad_input_pipe_300_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Zeropad_input_pipe_318_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Zeropad_input_pipe_336_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Zeropad_input_pipe_354_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Zeropad_input_pipe_372_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Zeropad_input_pipe_390_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Zeropad_input_pipe_408_inst_req_0;
      RPIPE_Zeropad_input_pipe_45_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_Zeropad_input_pipe_135_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_Zeropad_input_pipe_96_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_Zeropad_input_pipe_59_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_Zeropad_input_pipe_121_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_Zeropad_input_pipe_109_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_Zeropad_input_pipe_71_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Zeropad_input_pipe_84_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Zeropad_input_pipe_147_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Zeropad_input_pipe_160_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Zeropad_input_pipe_172_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Zeropad_input_pipe_185_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Zeropad_input_pipe_287_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Zeropad_input_pipe_300_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Zeropad_input_pipe_318_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Zeropad_input_pipe_336_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Zeropad_input_pipe_354_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Zeropad_input_pipe_372_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Zeropad_input_pipe_390_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Zeropad_input_pipe_408_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(19) <= RPIPE_Zeropad_input_pipe_45_inst_req_1;
      reqR_unguarded(18) <= RPIPE_Zeropad_input_pipe_135_inst_req_1;
      reqR_unguarded(17) <= RPIPE_Zeropad_input_pipe_96_inst_req_1;
      reqR_unguarded(16) <= RPIPE_Zeropad_input_pipe_59_inst_req_1;
      reqR_unguarded(15) <= RPIPE_Zeropad_input_pipe_121_inst_req_1;
      reqR_unguarded(14) <= RPIPE_Zeropad_input_pipe_109_inst_req_1;
      reqR_unguarded(13) <= RPIPE_Zeropad_input_pipe_71_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Zeropad_input_pipe_84_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Zeropad_input_pipe_147_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Zeropad_input_pipe_160_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Zeropad_input_pipe_172_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Zeropad_input_pipe_185_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Zeropad_input_pipe_287_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Zeropad_input_pipe_300_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Zeropad_input_pipe_318_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Zeropad_input_pipe_336_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Zeropad_input_pipe_354_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Zeropad_input_pipe_372_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Zeropad_input_pipe_390_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Zeropad_input_pipe_408_inst_req_1;
      RPIPE_Zeropad_input_pipe_45_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_Zeropad_input_pipe_135_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_Zeropad_input_pipe_96_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_Zeropad_input_pipe_59_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_Zeropad_input_pipe_121_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_Zeropad_input_pipe_109_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_Zeropad_input_pipe_71_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Zeropad_input_pipe_84_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Zeropad_input_pipe_147_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Zeropad_input_pipe_160_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Zeropad_input_pipe_172_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Zeropad_input_pipe_185_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Zeropad_input_pipe_287_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Zeropad_input_pipe_300_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Zeropad_input_pipe_318_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Zeropad_input_pipe_336_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Zeropad_input_pipe_354_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Zeropad_input_pipe_372_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Zeropad_input_pipe_390_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Zeropad_input_pipe_408_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      call_46 <= data_out(159 downto 152);
      call28_136 <= data_out(151 downto 144);
      call14_97 <= data_out(143 downto 136);
      call2_60 <= data_out(135 downto 128);
      call23_122 <= data_out(127 downto 120);
      call19_110 <= data_out(119 downto 112);
      call5_72 <= data_out(111 downto 104);
      call10_85 <= data_out(103 downto 96);
      call32_148 <= data_out(95 downto 88);
      call37_161 <= data_out(87 downto 80);
      call41_173 <= data_out(79 downto 72);
      call46_186 <= data_out(71 downto 64);
      call72_288 <= data_out(63 downto 56);
      call76_301 <= data_out(55 downto 48);
      call82_319 <= data_out(47 downto 40);
      call88_337 <= data_out(39 downto 32);
      call94_355 <= data_out(31 downto 24);
      call100_373 <= data_out(23 downto 16);
      call106_391 <= data_out(15 downto 8);
      call112_409 <= data_out(7 downto 0);
      Zeropad_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "Zeropad_input_pipe_read_0_gI", nreqs => 20, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Zeropad_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "Zeropad_input_pipe_read_0", data_width => 8,  num_reqs => 20,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Zeropad_input_pipe_pipe_read_req(0),
          oack => Zeropad_input_pipe_pipe_read_ack(0),
          odata => Zeropad_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Zeropad_output_pipe_1430_inst WPIPE_Zeropad_output_pipe_1433_inst WPIPE_Zeropad_output_pipe_1436_inst WPIPE_Zeropad_output_pipe_1439_inst WPIPE_Zeropad_output_pipe_1442_inst WPIPE_Zeropad_output_pipe_1445_inst WPIPE_Zeropad_output_pipe_1448_inst WPIPE_Zeropad_output_pipe_1451_inst WPIPE_Zeropad_output_pipe_1602_inst WPIPE_Zeropad_output_pipe_1605_inst WPIPE_Zeropad_output_pipe_1608_inst WPIPE_Zeropad_output_pipe_1611_inst WPIPE_Zeropad_output_pipe_1614_inst WPIPE_Zeropad_output_pipe_1617_inst WPIPE_Zeropad_output_pipe_1620_inst WPIPE_Zeropad_output_pipe_1623_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 15 downto 0);
      signal update_req, update_ack : BooleanArray( 15 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 15 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      sample_req_unguarded(15) <= WPIPE_Zeropad_output_pipe_1430_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_Zeropad_output_pipe_1433_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_Zeropad_output_pipe_1436_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Zeropad_output_pipe_1439_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Zeropad_output_pipe_1442_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Zeropad_output_pipe_1445_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Zeropad_output_pipe_1448_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Zeropad_output_pipe_1451_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Zeropad_output_pipe_1602_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Zeropad_output_pipe_1605_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Zeropad_output_pipe_1608_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Zeropad_output_pipe_1611_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Zeropad_output_pipe_1614_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Zeropad_output_pipe_1617_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Zeropad_output_pipe_1620_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Zeropad_output_pipe_1623_inst_req_0;
      WPIPE_Zeropad_output_pipe_1430_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_Zeropad_output_pipe_1433_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_Zeropad_output_pipe_1436_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Zeropad_output_pipe_1439_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Zeropad_output_pipe_1442_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Zeropad_output_pipe_1445_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Zeropad_output_pipe_1448_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Zeropad_output_pipe_1451_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Zeropad_output_pipe_1602_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Zeropad_output_pipe_1605_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Zeropad_output_pipe_1608_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Zeropad_output_pipe_1611_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Zeropad_output_pipe_1614_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Zeropad_output_pipe_1617_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Zeropad_output_pipe_1620_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Zeropad_output_pipe_1623_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(15) <= WPIPE_Zeropad_output_pipe_1430_inst_req_1;
      update_req_unguarded(14) <= WPIPE_Zeropad_output_pipe_1433_inst_req_1;
      update_req_unguarded(13) <= WPIPE_Zeropad_output_pipe_1436_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Zeropad_output_pipe_1439_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Zeropad_output_pipe_1442_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Zeropad_output_pipe_1445_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Zeropad_output_pipe_1448_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Zeropad_output_pipe_1451_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Zeropad_output_pipe_1602_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Zeropad_output_pipe_1605_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Zeropad_output_pipe_1608_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Zeropad_output_pipe_1611_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Zeropad_output_pipe_1614_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Zeropad_output_pipe_1617_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Zeropad_output_pipe_1620_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Zeropad_output_pipe_1623_inst_req_1;
      WPIPE_Zeropad_output_pipe_1430_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_Zeropad_output_pipe_1433_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_Zeropad_output_pipe_1436_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Zeropad_output_pipe_1439_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Zeropad_output_pipe_1442_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Zeropad_output_pipe_1445_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Zeropad_output_pipe_1448_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Zeropad_output_pipe_1451_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Zeropad_output_pipe_1602_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Zeropad_output_pipe_1605_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Zeropad_output_pipe_1608_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Zeropad_output_pipe_1611_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Zeropad_output_pipe_1614_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Zeropad_output_pipe_1617_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Zeropad_output_pipe_1620_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Zeropad_output_pipe_1623_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      data_in <= conv347_1429 & conv341_1419 & conv335_1409 & conv329_1399 & conv323_1389 & conv317_1379 & conv311_1369 & conv305_1359 & conv422_1601 & conv416_1591 & conv410_1581 & conv404_1571 & conv398_1561 & conv392_1551 & conv386_1541 & conv380_1531;
      Zeropad_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "Zeropad_output_pipe_write_0_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Zeropad_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "Zeropad_output_pipe", data_width => 8, num_reqs => 16, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Zeropad_output_pipe_pipe_write_req(0),
          oack => Zeropad_output_pipe_pipe_write_ack(0),
          odata => Zeropad_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_445_call call_stmt_1345_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_445_call_req_0;
      reqL_unguarded(0) <= call_stmt_1345_call_req_0;
      call_stmt_445_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1345_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_445_call_req_1;
      reqR_unguarded(0) <= call_stmt_1345_call_req_1;
      call_stmt_445_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1345_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call120_445 <= data_out(127 downto 64);
      call296_1345 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    Zeropad_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    Zeropad_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    Zeropad_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    Zeropad_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    Zeropad_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    Zeropad_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(14 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(14 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- declarations related to module zeropad
  component zeropad is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(14 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(14 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      Zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      Zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad
  signal zeropad_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad_start_req : std_logic;
  signal zeropad_start_ack : std_logic;
  signal zeropad_fin_req   : std_logic;
  signal zeropad_fin_ack : std_logic;
  -- aggregate signals for read from pipe Zeropad_input_pipe
  signal Zeropad_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal Zeropad_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal Zeropad_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Zeropad_output_pipe
  signal Zeropad_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal Zeropad_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal Zeropad_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(0 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(17 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(0 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(17 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  -- module zeropad
  zeropad_instance:zeropad-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad_start_req,
      start_ack => zeropad_start_ack,
      fin_req => zeropad_fin_req,
      fin_ack => zeropad_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(14 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(14 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      Zeropad_input_pipe_pipe_read_req => Zeropad_input_pipe_pipe_read_req(0 downto 0),
      Zeropad_input_pipe_pipe_read_ack => Zeropad_input_pipe_pipe_read_ack(0 downto 0),
      Zeropad_input_pipe_pipe_read_data => Zeropad_input_pipe_pipe_read_data(7 downto 0),
      Zeropad_output_pipe_pipe_write_req => Zeropad_output_pipe_pipe_write_req(0 downto 0),
      Zeropad_output_pipe_pipe_write_ack => Zeropad_output_pipe_pipe_write_ack(0 downto 0),
      Zeropad_output_pipe_pipe_write_data => Zeropad_output_pipe_pipe_write_data(7 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => zeropad_tag_in,
      tag_out => zeropad_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad_tag_in <= (others => '0');
  zeropad_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad_start_req, start_ack => zeropad_start_ack,  fin_req => zeropad_fin_req,  fin_ack => zeropad_fin_ack);
  Zeropad_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Zeropad_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => Zeropad_input_pipe_pipe_read_req,
      read_ack => Zeropad_input_pipe_pipe_read_ack,
      read_data => Zeropad_input_pipe_pipe_read_data,
      write_req => Zeropad_input_pipe_pipe_write_req,
      write_ack => Zeropad_input_pipe_pipe_write_ack,
      write_data => Zeropad_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Zeropad_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Zeropad_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => Zeropad_output_pipe_pipe_read_req,
      read_ack => Zeropad_output_pipe_pipe_read_ack,
      read_data => Zeropad_output_pipe_pipe_read_data,
      write_req => Zeropad_output_pipe_pipe_write_req,
      write_ack => Zeropad_output_pipe_pipe_write_ack,
      write_data => Zeropad_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 15,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 15,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
