-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package ahir_system_global_package is -- 
  constant KD1_1_base_address : std_logic_vector(13 downto 0) := "00000000000000";
  constant KD1_2_base_address : std_logic_vector(12 downto 0) := "0000000000000";
  constant KD2_1_base_address : std_logic_vector(15 downto 0) := "0000000000000000";
  constant KD2_2_base_address : std_logic_vector(14 downto 0) := "000000000000000";
  constant KD3_1_base_address : std_logic_vector(17 downto 0) := "000000000000000000";
  constant KD3_2_base_address : std_logic_vector(16 downto 0) := "00000000000000000";
  constant KE1_1_base_address : std_logic_vector(8 downto 0) := "000000000";
  constant KE1_2_base_address : std_logic_vector(12 downto 0) := "0000000000000";
  constant KE2_1_base_address : std_logic_vector(13 downto 0) := "00000000000000";
  constant KE2_2_base_address : std_logic_vector(14 downto 0) := "000000000000000";
  constant KE3_1_base_address : std_logic_vector(15 downto 0) := "0000000000000000";
  constant KE3_2_base_address : std_logic_vector(16 downto 0) := "00000000000000000";
  constant KL_base_address : std_logic_vector(8 downto 0) := "000000000";
  constant KM1_base_address : std_logic_vector(17 downto 0) := "000000000000000000";
  constant KM2_base_address : std_logic_vector(18 downto 0) := "0000000000000000000";
  constant KT1_base_address : std_logic_vector(13 downto 0) := "00000000000000";
  constant KT2_base_address : std_logic_vector(15 downto 0) := "0000000000000000";
  constant KT3_base_address : std_logic_vector(17 downto 0) := "000000000000000000";
  constant Tensor0_base_address : std_logic_vector(18 downto 0) := "0000000000000000000";
  constant Tensor1_base_address : std_logic_vector(19 downto 0) := "00000000000000000000";
  constant Tensor2_base_address : std_logic_vector(18 downto 0) := "0000000000000000000";
  constant Tensor3_base_address : std_logic_vector(17 downto 0) := "000000000000000000";
  constant Tensor4_base_address : std_logic_vector(16 downto 0) := "00000000000000000";
  -- 
end package ahir_system_global_package;
