-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity access_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    row_in : in  std_logic_vector(15 downto 0);
    chl_in : in  std_logic_vector(15 downto 0);
    ct : in  std_logic_vector(15 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    input_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
    input_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
    input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity access_T;
architecture access_T_arch of access_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 48)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal row_in_buffer :  std_logic_vector(15 downto 0);
  signal row_in_update_enable: Boolean;
  signal chl_in_buffer :  std_logic_vector(15 downto 0);
  signal chl_in_update_enable: Boolean;
  signal ct_buffer :  std_logic_vector(15 downto 0);
  signal ct_update_enable: Boolean;
  -- output port buffer signals
  signal access_T_CP_0_start: Boolean;
  signal access_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal W_fn3_330_delayed_13_0_359_inst_ack_1 : boolean;
  signal W_fn3_324_delayed_7_0_351_inst_req_1 : boolean;
  signal W_fetch_val3_332_delayed_13_0_362_inst_req_1 : boolean;
  signal W_fetch_val3_332_delayed_13_0_362_inst_ack_1 : boolean;
  signal addr_of_270_final_reg_ack_0 : boolean;
  signal W_fn3_330_delayed_13_0_359_inst_req_0 : boolean;
  signal W_fn3_330_delayed_13_0_359_inst_req_1 : boolean;
  signal W_fetch_val3_332_delayed_13_0_362_inst_req_0 : boolean;
  signal W_fetch_val3_332_delayed_13_0_362_inst_ack_0 : boolean;
  signal W_continue_307_delayed_1_0_323_inst_req_1 : boolean;
  signal ptr_deref_357_load_0_req_1 : boolean;
  signal W_fn2_257_delayed_7_0_272_inst_ack_1 : boolean;
  signal W_fn2_257_delayed_7_0_272_inst_req_1 : boolean;
  signal ptr_deref_49_load_0_req_0 : boolean;
  signal ptr_deref_49_load_0_ack_0 : boolean;
  signal addr_of_270_final_reg_req_0 : boolean;
  signal ptr_deref_49_load_0_req_1 : boolean;
  signal ptr_deref_49_load_0_ack_1 : boolean;
  signal WPIPE_input_pipe2_292_inst_ack_1 : boolean;
  signal WPIPE_input_pipe2_292_inst_req_1 : boolean;
  signal array_obj_ref_58_index_offset_req_0 : boolean;
  signal array_obj_ref_58_index_offset_ack_0 : boolean;
  signal array_obj_ref_58_index_offset_req_1 : boolean;
  signal array_obj_ref_58_index_offset_ack_1 : boolean;
  signal addr_of_349_final_reg_ack_0 : boolean;
  signal addr_of_349_final_reg_req_0 : boolean;
  signal addr_of_59_final_reg_req_0 : boolean;
  signal addr_of_59_final_reg_ack_0 : boolean;
  signal W_fn2_263_delayed_13_0_280_inst_ack_0 : boolean;
  signal addr_of_59_final_reg_req_1 : boolean;
  signal addr_of_59_final_reg_ack_1 : boolean;
  signal WPIPE_input_pipe2_292_inst_ack_0 : boolean;
  signal W_fn2_257_delayed_7_0_272_inst_ack_0 : boolean;
  signal W_fn2_257_delayed_7_0_272_inst_req_0 : boolean;
  signal ptr_deref_63_load_0_req_0 : boolean;
  signal ptr_deref_63_load_0_ack_0 : boolean;
  signal W_fn2_263_delayed_13_0_280_inst_req_0 : boolean;
  signal ptr_deref_63_load_0_req_1 : boolean;
  signal ptr_deref_63_load_0_ack_1 : boolean;
  signal WPIPE_input_pipe2_292_inst_req_0 : boolean;
  signal W_fn3_324_delayed_7_0_351_inst_ack_0 : boolean;
  signal array_obj_ref_72_index_offset_req_0 : boolean;
  signal array_obj_ref_72_index_offset_ack_0 : boolean;
  signal array_obj_ref_72_index_offset_req_1 : boolean;
  signal array_obj_ref_72_index_offset_ack_1 : boolean;
  signal type_cast_90_inst_req_0 : boolean;
  signal type_cast_90_inst_ack_0 : boolean;
  signal type_cast_90_inst_req_1 : boolean;
  signal type_cast_90_inst_ack_1 : boolean;
  signal addr_of_73_final_reg_req_0 : boolean;
  signal addr_of_73_final_reg_ack_0 : boolean;
  signal addr_of_73_final_reg_req_1 : boolean;
  signal addr_of_73_final_reg_ack_1 : boolean;
  signal ptr_deref_77_load_0_req_0 : boolean;
  signal ptr_deref_77_load_0_ack_0 : boolean;
  signal ptr_deref_77_load_0_req_1 : boolean;
  signal ptr_deref_77_load_0_ack_1 : boolean;
  signal ptr_deref_357_load_0_ack_0 : boolean;
  signal W_continue_307_delayed_1_0_323_inst_ack_0 : boolean;
  signal do_while_stmt_79_branch_req_0 : boolean;
  signal array_obj_ref_269_index_offset_ack_1 : boolean;
  signal W_continue_307_delayed_1_0_323_inst_req_0 : boolean;
  signal W_fn3_324_delayed_7_0_351_inst_req_0 : boolean;
  signal phi_stmt_81_req_0 : boolean;
  signal phi_stmt_81_req_1 : boolean;
  signal array_obj_ref_269_index_offset_req_1 : boolean;
  signal phi_stmt_81_ack_0 : boolean;
  signal n_address1_174_83_buf_req_0 : boolean;
  signal n_address1_174_83_buf_ack_0 : boolean;
  signal n_address1_174_83_buf_req_1 : boolean;
  signal n_address1_174_83_buf_ack_1 : boolean;
  signal addr_of_270_final_reg_ack_1 : boolean;
  signal phi_stmt_86_req_0 : boolean;
  signal phi_stmt_86_req_1 : boolean;
  signal array_obj_ref_269_index_offset_ack_0 : boolean;
  signal phi_stmt_86_ack_0 : boolean;
  signal addr_of_270_final_reg_req_1 : boolean;
  signal n_address2_248_88_buf_req_0 : boolean;
  signal n_address2_248_88_buf_ack_0 : boolean;
  signal array_obj_ref_269_index_offset_req_0 : boolean;
  signal n_address2_248_88_buf_req_1 : boolean;
  signal n_address2_248_88_buf_ack_1 : boolean;
  signal phi_stmt_113_req_0 : boolean;
  signal phi_stmt_113_req_1 : boolean;
  signal phi_stmt_113_ack_0 : boolean;
  signal ptr_deref_357_load_0_req_0 : boolean;
  signal ptr_deref_278_load_0_ack_1 : boolean;
  signal ptr_deref_278_load_0_req_1 : boolean;
  signal phi_stmt_91_req_0 : boolean;
  signal phi_stmt_91_req_1 : boolean;
  signal phi_stmt_91_ack_0 : boolean;
  signal n_address3_322_93_buf_req_0 : boolean;
  signal n_address3_322_93_buf_ack_0 : boolean;
  signal n_address3_322_93_buf_req_1 : boolean;
  signal n_address3_322_93_buf_ack_1 : boolean;
  signal type_cast_95_inst_req_0 : boolean;
  signal type_cast_95_inst_ack_0 : boolean;
  signal type_cast_95_inst_req_1 : boolean;
  signal type_cast_95_inst_ack_1 : boolean;
  signal addr_of_349_final_reg_ack_1 : boolean;
  signal addr_of_349_final_reg_req_1 : boolean;
  signal W_fn3_330_delayed_13_0_359_inst_ack_0 : boolean;
  signal phi_stmt_96_req_0 : boolean;
  signal phi_stmt_96_req_1 : boolean;
  signal phi_stmt_96_ack_0 : boolean;
  signal W_fetch_val2_265_delayed_13_0_283_inst_ack_1 : boolean;
  signal W_fetch_val2_265_delayed_13_0_283_inst_req_1 : boolean;
  signal n_mycounter_141_98_buf_req_0 : boolean;
  signal n_mycounter_141_98_buf_ack_0 : boolean;
  signal ptr_deref_357_load_0_ack_1 : boolean;
  signal n_mycounter_141_98_buf_req_1 : boolean;
  signal n_mycounter_141_98_buf_ack_1 : boolean;
  signal W_fn3_324_delayed_7_0_351_inst_ack_1 : boolean;
  signal W_fetch_val2_265_delayed_13_0_283_inst_ack_0 : boolean;
  signal W_fetch_val2_265_delayed_13_0_283_inst_req_0 : boolean;
  signal ptr_deref_278_load_0_ack_0 : boolean;
  signal ptr_deref_278_load_0_req_0 : boolean;
  signal array_obj_ref_348_index_offset_ack_1 : boolean;
  signal array_obj_ref_348_index_offset_req_1 : boolean;
  signal phi_stmt_101_req_0 : boolean;
  signal phi_stmt_101_req_1 : boolean;
  signal array_obj_ref_348_index_offset_ack_0 : boolean;
  signal phi_stmt_101_ack_0 : boolean;
  signal n_fetch_val1_217_103_buf_req_0 : boolean;
  signal W_fn2_263_delayed_13_0_280_inst_ack_1 : boolean;
  signal n_fetch_val1_217_103_buf_ack_0 : boolean;
  signal n_fetch_val1_217_103_buf_req_1 : boolean;
  signal n_fetch_val1_217_103_buf_ack_1 : boolean;
  signal array_obj_ref_348_index_offset_req_0 : boolean;
  signal my_fetch1_50_104_buf_req_0 : boolean;
  signal W_fn2_263_delayed_13_0_280_inst_req_1 : boolean;
  signal my_fetch1_50_104_buf_ack_0 : boolean;
  signal W_continue_307_delayed_1_0_323_inst_ack_1 : boolean;
  signal my_fetch1_50_104_buf_req_1 : boolean;
  signal my_fetch1_50_104_buf_ack_1 : boolean;
  signal phi_stmt_105_req_0 : boolean;
  signal phi_stmt_105_req_1 : boolean;
  signal phi_stmt_105_ack_0 : boolean;
  signal n_fetch_val2_291_107_buf_req_0 : boolean;
  signal n_fetch_val2_291_107_buf_ack_0 : boolean;
  signal n_fetch_val2_291_107_buf_req_1 : boolean;
  signal n_fetch_val2_291_107_buf_ack_1 : boolean;
  signal my_fetch2_64_108_buf_req_0 : boolean;
  signal my_fetch2_64_108_buf_ack_0 : boolean;
  signal my_fetch2_64_108_buf_req_1 : boolean;
  signal my_fetch2_64_108_buf_ack_1 : boolean;
  signal phi_stmt_109_req_0 : boolean;
  signal phi_stmt_109_req_1 : boolean;
  signal phi_stmt_109_ack_0 : boolean;
  signal n_fetch_val3_370_111_buf_req_0 : boolean;
  signal n_fetch_val3_370_111_buf_ack_0 : boolean;
  signal n_fetch_val3_370_111_buf_req_1 : boolean;
  signal n_fetch_val3_370_111_buf_ack_1 : boolean;
  signal my_fetch3_78_112_buf_req_0 : boolean;
  signal my_fetch3_78_112_buf_ack_0 : boolean;
  signal my_fetch3_78_112_buf_req_1 : boolean;
  signal my_fetch3_78_112_buf_ack_1 : boolean;
  signal n_row1_169_115_buf_req_0 : boolean;
  signal n_row1_169_115_buf_ack_0 : boolean;
  signal n_row1_169_115_buf_req_1 : boolean;
  signal n_row1_169_115_buf_ack_1 : boolean;
  signal phi_stmt_118_req_1 : boolean;
  signal phi_stmt_118_req_0 : boolean;
  signal phi_stmt_118_ack_0 : boolean;
  signal n_row2_243_122_buf_req_0 : boolean;
  signal n_row2_243_122_buf_ack_0 : boolean;
  signal n_row2_243_122_buf_req_1 : boolean;
  signal n_row2_243_122_buf_ack_1 : boolean;
  signal phi_stmt_123_req_1 : boolean;
  signal phi_stmt_123_req_0 : boolean;
  signal phi_stmt_123_ack_0 : boolean;
  signal n_row3_317_127_buf_req_0 : boolean;
  signal n_row3_317_127_buf_ack_0 : boolean;
  signal n_row3_317_127_buf_req_1 : boolean;
  signal n_row3_317_127_buf_ack_1 : boolean;
  signal W_continue_183_delayed_1_0_175_inst_req_0 : boolean;
  signal W_continue_183_delayed_1_0_175_inst_ack_0 : boolean;
  signal W_continue_183_delayed_1_0_175_inst_req_1 : boolean;
  signal W_continue_183_delayed_1_0_175_inst_ack_1 : boolean;
  signal array_obj_ref_195_index_offset_req_0 : boolean;
  signal array_obj_ref_195_index_offset_ack_0 : boolean;
  signal array_obj_ref_195_index_offset_req_1 : boolean;
  signal array_obj_ref_195_index_offset_ack_1 : boolean;
  signal addr_of_196_final_reg_req_0 : boolean;
  signal addr_of_196_final_reg_ack_0 : boolean;
  signal addr_of_196_final_reg_req_1 : boolean;
  signal addr_of_196_final_reg_ack_1 : boolean;
  signal W_fn1_195_delayed_7_0_198_inst_req_0 : boolean;
  signal W_fn1_195_delayed_7_0_198_inst_ack_0 : boolean;
  signal W_fn1_195_delayed_7_0_198_inst_req_1 : boolean;
  signal W_fn1_195_delayed_7_0_198_inst_ack_1 : boolean;
  signal ptr_deref_204_load_0_req_0 : boolean;
  signal ptr_deref_204_load_0_ack_0 : boolean;
  signal ptr_deref_204_load_0_req_1 : boolean;
  signal ptr_deref_204_load_0_ack_1 : boolean;
  signal W_fn1_201_delayed_13_0_206_inst_req_0 : boolean;
  signal W_fn1_201_delayed_13_0_206_inst_ack_0 : boolean;
  signal W_fn1_201_delayed_13_0_206_inst_req_1 : boolean;
  signal W_fn1_201_delayed_13_0_206_inst_ack_1 : boolean;
  signal W_fetch_val1_203_delayed_13_0_209_inst_req_0 : boolean;
  signal W_fetch_val1_203_delayed_13_0_209_inst_ack_0 : boolean;
  signal W_fetch_val1_203_delayed_13_0_209_inst_req_1 : boolean;
  signal W_fetch_val1_203_delayed_13_0_209_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_218_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_218_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_218_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_218_inst_ack_1 : boolean;
  signal W_continue_245_delayed_1_0_249_inst_req_0 : boolean;
  signal W_continue_245_delayed_1_0_249_inst_ack_0 : boolean;
  signal W_continue_245_delayed_1_0_249_inst_req_1 : boolean;
  signal W_continue_245_delayed_1_0_249_inst_ack_1 : boolean;
  signal WPIPE_input_pipe3_372_inst_req_0 : boolean;
  signal WPIPE_input_pipe3_372_inst_ack_0 : boolean;
  signal WPIPE_input_pipe3_372_inst_req_1 : boolean;
  signal WPIPE_input_pipe3_372_inst_ack_1 : boolean;
  signal do_while_stmt_79_branch_ack_0 : boolean;
  signal do_while_stmt_79_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "access_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 48) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(15 downto 0) <= row_in;
  row_in_buffer <= in_buffer_data_out(15 downto 0);
  in_buffer_data_in(31 downto 16) <= chl_in;
  chl_in_buffer <= in_buffer_data_out(31 downto 16);
  in_buffer_data_in(47 downto 32) <= ct;
  ct_buffer <= in_buffer_data_out(47 downto 32);
  in_buffer_data_in(tag_length + 47 downto 48) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 47 downto 48);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  access_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "access_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  access_T_CP_0: Block -- control-path 
    signal access_T_CP_0_elements: BooleanArray(316 downto 0);
    -- 
  begin -- 
    access_T_CP_0_elements(0) <= access_T_CP_0_start;
    access_T_CP_0_symbol <= access_T_CP_0_elements(1);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	10 
    -- CP-element group 0: 	11 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	15 
    -- CP-element group 0:  members (79) 
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_index_scale_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_index_scale_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_26/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/branch_block_stmt_26__entry__
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78__entry__
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_59_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_index_resized_1
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_index_scaled_1
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_index_computed_1
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_index_resize_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_index_resize_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_index_resize_1/index_resize_req
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_final_index_sum_regn_update_start
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_59_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_59_complete/req
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_73_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_index_resized_1
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_index_scaled_1
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_index_computed_1
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_index_resize_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_index_resize_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_index_resize_1/index_resize_req
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_index_scale_1/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_index_scale_1/$exit
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_final_index_sum_regn_update_start
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_73_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_73_complete/req
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_update_start_
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Update/word_access_complete/word_0/cr
      -- 
    rr_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => ptr_deref_49_load_0_req_0); -- 
    cr_58_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_58_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => ptr_deref_49_load_0_req_1); -- 
    req_89_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_89_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_58_index_offset_req_0); -- 
    req_94_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_94_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_58_index_offset_req_1); -- 
    req_109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => addr_of_59_final_reg_req_1); -- 
    cr_154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => ptr_deref_63_load_0_req_1); -- 
    req_185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_72_index_offset_req_0); -- 
    req_190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => array_obj_ref_72_index_offset_req_1); -- 
    req_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => addr_of_73_final_reg_req_1); -- 
    cr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(0), ack => ptr_deref_77_load_0_req_1); -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	316 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_26/$exit
      -- CP-element group 1: 	 branch_block_stmt_26/branch_block_stmt_26__exit__
      -- CP-element group 1: 	 branch_block_stmt_26/do_while_stmt_79__exit__
      -- 
    access_T_CP_0_elements(1) <= access_T_CP_0_elements(316);
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Sample/word_access_start/$exit
      -- CP-element group 2: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Sample/word_access_start/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Sample/word_access_start/word_0/ra
      -- 
    ra_48_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_49_load_0_ack_0, ack => access_T_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	16 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Update/word_access_complete/$exit
      -- CP-element group 3: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Update/word_access_complete/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Update/word_access_complete/word_0/ca
      -- CP-element group 3: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Update/ptr_deref_49_Merge/$entry
      -- CP-element group 3: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Update/ptr_deref_49_Merge/$exit
      -- CP-element group 3: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Update/ptr_deref_49_Merge/merge_req
      -- CP-element group 3: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_49_Update/ptr_deref_49_Merge/merge_ack
      -- 
    ca_59_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_49_load_0_ack_1, ack => access_T_CP_0_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	16 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_final_index_sum_regn_sample_complete
      -- CP-element group 4: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_final_index_sum_regn_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_final_index_sum_regn_Sample/ack
      -- 
    ack_90_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_58_index_offset_ack_0, ack => access_T_CP_0_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (11) 
      -- CP-element group 5: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_59_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_root_address_calculated
      -- CP-element group 5: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_offset_calculated
      -- CP-element group 5: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_final_index_sum_regn_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_final_index_sum_regn_Update/ack
      -- CP-element group 5: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_base_plus_offset/$entry
      -- CP-element group 5: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_base_plus_offset/$exit
      -- CP-element group 5: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_base_plus_offset/sum_rename_req
      -- CP-element group 5: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_58_base_plus_offset/sum_rename_ack
      -- CP-element group 5: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_59_request/$entry
      -- CP-element group 5: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_59_request/req
      -- 
    ack_95_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_58_index_offset_ack_1, ack => access_T_CP_0_elements(5)); -- 
    req_104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(5), ack => addr_of_59_final_reg_req_0); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_59_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_59_request/$exit
      -- CP-element group 6: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_59_request/ack
      -- 
    ack_105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_59_final_reg_ack_0, ack => access_T_CP_0_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (24) 
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_59_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_59_complete/$exit
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_59_complete/ack
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_base_address_calculated
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_word_address_calculated
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_root_address_calculated
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_base_address_resized
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_base_addr_resize/$entry
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_base_addr_resize/$exit
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_base_addr_resize/base_resize_req
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_base_addr_resize/base_resize_ack
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_base_plus_offset/$entry
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_base_plus_offset/$exit
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_base_plus_offset/sum_rename_req
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_base_plus_offset/sum_rename_ack
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_word_addrgen/$entry
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_word_addrgen/$exit
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_word_addrgen/root_register_req
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_word_addrgen/root_register_ack
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Sample/word_access_start/$entry
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Sample/word_access_start/word_0/$entry
      -- CP-element group 7: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Sample/word_access_start/word_0/rr
      -- 
    ack_110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_59_final_reg_ack_1, ack => access_T_CP_0_elements(7)); -- 
    rr_143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(7), ack => ptr_deref_63_load_0_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (5) 
      -- CP-element group 8: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Sample/word_access_start/$exit
      -- CP-element group 8: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Sample/word_access_start/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Sample/word_access_start/word_0/ra
      -- 
    ra_144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_63_load_0_ack_0, ack => access_T_CP_0_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	16 
    -- CP-element group 9:  members (9) 
      -- CP-element group 9: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Update/word_access_complete/$exit
      -- CP-element group 9: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Update/word_access_complete/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Update/word_access_complete/word_0/ca
      -- CP-element group 9: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Update/ptr_deref_63_Merge/$entry
      -- CP-element group 9: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Update/ptr_deref_63_Merge/$exit
      -- CP-element group 9: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Update/ptr_deref_63_Merge/merge_req
      -- CP-element group 9: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_63_Update/ptr_deref_63_Merge/merge_ack
      -- 
    ca_155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_63_load_0_ack_1, ack => access_T_CP_0_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	16 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_final_index_sum_regn_sample_complete
      -- CP-element group 10: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_final_index_sum_regn_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_final_index_sum_regn_Sample/ack
      -- 
    ack_186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_72_index_offset_ack_0, ack => access_T_CP_0_elements(10)); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (11) 
      -- CP-element group 11: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_base_plus_offset/$entry
      -- CP-element group 11: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_base_plus_offset/$exit
      -- CP-element group 11: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_base_plus_offset/sum_rename_req
      -- CP-element group 11: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_base_plus_offset/sum_rename_ack
      -- CP-element group 11: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_73_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_root_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_offset_calculated
      -- CP-element group 11: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_final_index_sum_regn_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/array_obj_ref_72_final_index_sum_regn_Update/ack
      -- CP-element group 11: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_73_request/$entry
      -- CP-element group 11: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_73_request/req
      -- 
    ack_191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_72_index_offset_ack_1, ack => access_T_CP_0_elements(11)); -- 
    req_200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(11), ack => addr_of_73_final_reg_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_73_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_73_request/$exit
      -- CP-element group 12: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_73_request/ack
      -- 
    ack_201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_73_final_reg_ack_0, ack => access_T_CP_0_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (24) 
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_73_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_73_complete/$exit
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/addr_of_73_complete/ack
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_base_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_word_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_root_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_base_address_resized
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_base_addr_resize/$entry
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_base_addr_resize/$exit
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_base_addr_resize/base_resize_req
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_base_addr_resize/base_resize_ack
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_base_plus_offset/$entry
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_base_plus_offset/$exit
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_base_plus_offset/sum_rename_req
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_base_plus_offset/sum_rename_ack
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_word_addrgen/$entry
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_word_addrgen/$exit
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_word_addrgen/root_register_req
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_word_addrgen/root_register_ack
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Sample/word_access_start/$entry
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Sample/word_access_start/word_0/$entry
      -- CP-element group 13: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Sample/word_access_start/word_0/rr
      -- 
    ack_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_73_final_reg_ack_1, ack => access_T_CP_0_elements(13)); -- 
    rr_239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(13), ack => ptr_deref_77_load_0_req_0); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Sample/word_access_start/$exit
      -- CP-element group 14: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Sample/word_access_start/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Sample/word_access_start/word_0/ra
      -- 
    ra_240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_77_load_0_ack_0, ack => access_T_CP_0_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	0 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Update/word_access_complete/$exit
      -- CP-element group 15: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Update/word_access_complete/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Update/word_access_complete/word_0/ca
      -- CP-element group 15: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Update/ptr_deref_77_Merge/$entry
      -- CP-element group 15: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Update/ptr_deref_77_Merge/$exit
      -- CP-element group 15: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Update/ptr_deref_77_Merge/merge_req
      -- CP-element group 15: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/ptr_deref_77_Update/ptr_deref_77_Merge/merge_ack
      -- 
    ca_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_77_load_0_ack_1, ack => access_T_CP_0_elements(15)); -- 
    -- CP-element group 16:  join  transition  place  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	3 
    -- CP-element group 16: 	4 
    -- CP-element group 16: 	9 
    -- CP-element group 16: 	10 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78__exit__
      -- CP-element group 16: 	 branch_block_stmt_26/do_while_stmt_79__entry__
      -- CP-element group 16: 	 branch_block_stmt_26/assign_stmt_33_to_assign_stmt_78/$exit
      -- 
    access_T_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(3) & access_T_CP_0_elements(4) & access_T_CP_0_elements(9) & access_T_CP_0_elements(10) & access_T_CP_0_elements(15);
      gj_access_T_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  transition  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	23 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_26/do_while_stmt_79/$entry
      -- CP-element group 17: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79__entry__
      -- 
    access_T_CP_0_elements(17) <= access_T_CP_0_elements(16);
    -- CP-element group 18:  merge  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	316 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79__exit__
      -- 
    -- Element group access_T_CP_0_elements(18) is bound as output of CP function.
    -- CP-element group 19:  merge  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_26/do_while_stmt_79/loop_back
      -- 
    -- Element group access_T_CP_0_elements(19) is bound as output of CP function.
    -- CP-element group 20:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	25 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	314 
    -- CP-element group 20: 	315 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_79/condition_done
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_79/loop_exit/$entry
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_79/loop_taken/$entry
      -- 
    access_T_CP_0_elements(20) <= access_T_CP_0_elements(25);
    -- CP-element group 21:  branch  place  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	313 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_26/do_while_stmt_79/loop_body_done
      -- 
    access_T_CP_0_elements(21) <= access_T_CP_0_elements(313);
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	95 
    -- CP-element group 22: 	114 
    -- CP-element group 22: 	76 
    -- CP-element group 22: 	55 
    -- CP-element group 22: 	36 
    -- CP-element group 22: 	133 
    -- CP-element group 22: 	152 
    -- CP-element group 22: 	171 
    -- CP-element group 22: 	190 
    -- CP-element group 22: 	209 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/back_edge_to_loop_body
      -- 
    access_T_CP_0_elements(22) <= access_T_CP_0_elements(19);
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	17 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	97 
    -- CP-element group 23: 	116 
    -- CP-element group 23: 	78 
    -- CP-element group 23: 	57 
    -- CP-element group 23: 	38 
    -- CP-element group 23: 	135 
    -- CP-element group 23: 	154 
    -- CP-element group 23: 	173 
    -- CP-element group 23: 	192 
    -- CP-element group 23: 	211 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/first_time_through_loop_body
      -- 
    access_T_CP_0_elements(23) <= access_T_CP_0_elements(17);
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	91 
    -- CP-element group 24: 	92 
    -- CP-element group 24: 	108 
    -- CP-element group 24: 	109 
    -- CP-element group 24: 	71 
    -- CP-element group 24: 	50 
    -- CP-element group 24: 	70 
    -- CP-element group 24: 	49 
    -- CP-element group 24: 	30 
    -- CP-element group 24: 	31 
    -- CP-element group 24: 	127 
    -- CP-element group 24: 	128 
    -- CP-element group 24: 	146 
    -- CP-element group 24: 	147 
    -- CP-element group 24: 	165 
    -- CP-element group 24: 	166 
    -- CP-element group 24: 	184 
    -- CP-element group 24: 	185 
    -- CP-element group 24: 	203 
    -- CP-element group 24: 	204 
    -- CP-element group 24: 	227 
    -- CP-element group 24: 	228 
    -- CP-element group 24: 	257 
    -- CP-element group 24: 	258 
    -- CP-element group 24: 	287 
    -- CP-element group 24: 	288 
    -- CP-element group 24: 	312 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/$entry
      -- CP-element group 24: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/loop_body_start
      -- 
    -- Element group access_T_CP_0_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	94 
    -- CP-element group 25: 	29 
    -- CP-element group 25: 	170 
    -- CP-element group 25: 	312 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	20 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/condition_evaluated
      -- 
    condition_evaluated_271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(25), ack => do_while_stmt_79_branch_req_0); -- 
    access_T_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(94) & access_T_CP_0_elements(29) & access_T_CP_0_elements(170) & access_T_CP_0_elements(312);
      gj_access_T_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	91 
    -- CP-element group 26: 	108 
    -- CP-element group 26: 	70 
    -- CP-element group 26: 	49 
    -- CP-element group 26: 	30 
    -- CP-element group 26: 	127 
    -- CP-element group 26: 	146 
    -- CP-element group 26: 	165 
    -- CP-element group 26: 	184 
    -- CP-element group 26: 	203 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	29 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	110 
    -- CP-element group 26: 	51 
    -- CP-element group 26: 	72 
    -- CP-element group 26: 	32 
    -- CP-element group 26: 	129 
    -- CP-element group 26: 	148 
    -- CP-element group 26: 	167 
    -- CP-element group 26: 	186 
    -- CP-element group 26: 	205 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/aggregated_phi_sample_req
      -- CP-element group 26: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_96_sample_start__ps
      -- 
    access_T_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 1);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= access_T_CP_0_elements(91) & access_T_CP_0_elements(108) & access_T_CP_0_elements(70) & access_T_CP_0_elements(49) & access_T_CP_0_elements(30) & access_T_CP_0_elements(127) & access_T_CP_0_elements(146) & access_T_CP_0_elements(165) & access_T_CP_0_elements(184) & access_T_CP_0_elements(203) & access_T_CP_0_elements(29);
      gj_access_T_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	93 
    -- CP-element group 27: 	111 
    -- CP-element group 27: 	73 
    -- CP-element group 27: 	52 
    -- CP-element group 27: 	33 
    -- CP-element group 27: 	130 
    -- CP-element group 27: 	149 
    -- CP-element group 27: 	168 
    -- CP-element group 27: 	187 
    -- CP-element group 27: 	206 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	238 
    -- CP-element group 27: 	242 
    -- CP-element group 27: 	246 
    -- CP-element group 27: 	268 
    -- CP-element group 27: 	272 
    -- CP-element group 27: 	276 
    -- CP-element group 27: 	298 
    -- CP-element group 27: 	302 
    -- CP-element group 27: 	306 
    -- CP-element group 27: 	313 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	91 
    -- CP-element group 27: 	108 
    -- CP-element group 27: 	70 
    -- CP-element group 27: 	49 
    -- CP-element group 27: 	30 
    -- CP-element group 27: 	127 
    -- CP-element group 27: 	146 
    -- CP-element group 27: 	165 
    -- CP-element group 27: 	184 
    -- CP-element group 27: 	203 
    -- CP-element group 27:  members (11) 
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/aggregated_phi_sample_ack
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_81_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_86_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_91_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_96_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_101_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_105_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_109_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_113_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_118_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_123_sample_completed_
      -- 
    access_T_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= access_T_CP_0_elements(93) & access_T_CP_0_elements(111) & access_T_CP_0_elements(73) & access_T_CP_0_elements(52) & access_T_CP_0_elements(33) & access_T_CP_0_elements(130) & access_T_CP_0_elements(149) & access_T_CP_0_elements(168) & access_T_CP_0_elements(187) & access_T_CP_0_elements(206);
      gj_access_T_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	92 
    -- CP-element group 28: 	109 
    -- CP-element group 28: 	71 
    -- CP-element group 28: 	50 
    -- CP-element group 28: 	31 
    -- CP-element group 28: 	128 
    -- CP-element group 28: 	147 
    -- CP-element group 28: 	166 
    -- CP-element group 28: 	185 
    -- CP-element group 28: 	204 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	112 
    -- CP-element group 28: 	74 
    -- CP-element group 28: 	53 
    -- CP-element group 28: 	34 
    -- CP-element group 28: 	131 
    -- CP-element group 28: 	150 
    -- CP-element group 28: 	169 
    -- CP-element group 28: 	188 
    -- CP-element group 28: 	207 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/aggregated_phi_update_req
      -- CP-element group 28: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_96_update_start__ps
      -- 
    access_T_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= access_T_CP_0_elements(92) & access_T_CP_0_elements(109) & access_T_CP_0_elements(71) & access_T_CP_0_elements(50) & access_T_CP_0_elements(31) & access_T_CP_0_elements(128) & access_T_CP_0_elements(147) & access_T_CP_0_elements(166) & access_T_CP_0_elements(185) & access_T_CP_0_elements(204);
      gj_access_T_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	94 
    -- CP-element group 29: 	113 
    -- CP-element group 29: 	75 
    -- CP-element group 29: 	54 
    -- CP-element group 29: 	35 
    -- CP-element group 29: 	132 
    -- CP-element group 29: 	151 
    -- CP-element group 29: 	170 
    -- CP-element group 29: 	189 
    -- CP-element group 29: 	208 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	25 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	26 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/aggregated_phi_update_ack
      -- 
    access_T_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= access_T_CP_0_elements(94) & access_T_CP_0_elements(113) & access_T_CP_0_elements(75) & access_T_CP_0_elements(54) & access_T_CP_0_elements(35) & access_T_CP_0_elements(132) & access_T_CP_0_elements(151) & access_T_CP_0_elements(170) & access_T_CP_0_elements(189) & access_T_CP_0_elements(208);
      gj_access_T_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	24 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	26 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_81_sample_start_
      -- 
    access_T_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27);
      gj_access_T_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	24 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	35 
    -- CP-element group 31: 	229 
    -- CP-element group 31: 	235 
    -- CP-element group 31: 	243 
    -- CP-element group 31: 	250 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	28 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_81_update_start_
      -- 
    access_T_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(35) & access_T_CP_0_elements(229) & access_T_CP_0_elements(235) & access_T_CP_0_elements(243) & access_T_CP_0_elements(250);
      gj_access_T_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	26 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_81_sample_start__ps
      -- 
    access_T_CP_0_elements(32) <= access_T_CP_0_elements(26);
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	27 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_81_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(33) is bound as output of CP function.
    -- CP-element group 34:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	28 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_81_update_start__ps
      -- 
    access_T_CP_0_elements(34) <= access_T_CP_0_elements(28);
    -- CP-element group 35:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	29 
    -- CP-element group 35: 	229 
    -- CP-element group 35: 	233 
    -- CP-element group 35: 	241 
    -- CP-element group 35: 	249 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	31 
    -- CP-element group 35:  members (15) 
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_81_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_81_update_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_index_resized_1
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_index_scaled_1
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_index_computed_1
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_index_resize_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_index_resize_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_index_resize_1/index_resize_req
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_index_resize_1/index_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_index_scale_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_index_scale_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_index_scale_1/scale_rename_req
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_index_scale_1/scale_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_final_index_sum_regn_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_final_index_sum_regn_Sample/req
      -- 
    req_805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(35), ack => array_obj_ref_195_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(35) is bound as output of CP function.
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	22 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_81_loopback_trigger
      -- 
    access_T_CP_0_elements(36) <= access_T_CP_0_elements(22);
    -- CP-element group 37:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_81_loopback_sample_req
      -- CP-element group 37: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_81_loopback_sample_req_ps
      -- 
    phi_stmt_81_loopback_sample_req_286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_81_loopback_sample_req_286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(37), ack => phi_stmt_81_req_0); -- 
    -- Element group access_T_CP_0_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	23 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_81_entry_trigger
      -- 
    access_T_CP_0_elements(38) <= access_T_CP_0_elements(23);
    -- CP-element group 39:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_81_entry_sample_req
      -- CP-element group 39: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_81_entry_sample_req_ps
      -- 
    phi_stmt_81_entry_sample_req_289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_81_entry_sample_req_289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(39), ack => phi_stmt_81_req_1); -- 
    -- Element group access_T_CP_0_elements(39) is bound as output of CP function.
    -- CP-element group 40:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (2) 
      -- CP-element group 40: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_81_phi_mux_ack
      -- CP-element group 40: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_81_phi_mux_ack_ps
      -- 
    phi_stmt_81_phi_mux_ack_292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_81_ack_0, ack => access_T_CP_0_elements(40)); -- 
    -- CP-element group 41:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (4) 
      -- CP-element group 41: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address1_83_sample_start__ps
      -- CP-element group 41: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address1_83_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address1_83_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address1_83_Sample/req
      -- 
    req_305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(41), ack => n_address1_174_83_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (4) 
      -- CP-element group 42: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address1_83_update_start__ps
      -- CP-element group 42: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address1_83_update_start_
      -- CP-element group 42: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address1_83_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address1_83_Update/req
      -- 
    req_310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(42), ack => n_address1_174_83_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(42) is bound as output of CP function.
    -- CP-element group 43:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address1_83_sample_completed__ps
      -- CP-element group 43: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address1_83_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address1_83_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address1_83_Sample/ack
      -- 
    ack_306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_174_83_buf_ack_0, ack => access_T_CP_0_elements(43)); -- 
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (4) 
      -- CP-element group 44: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address1_83_update_completed__ps
      -- CP-element group 44: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address1_83_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address1_83_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address1_83_Update/ack
      -- 
    ack_311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_174_83_buf_ack_1, ack => access_T_CP_0_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_85_sample_start__ps
      -- CP-element group 45: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_85_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_85_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_85_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_85_update_start__ps
      -- CP-element group 46: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_85_update_start_
      -- 
    -- Element group access_T_CP_0_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_85_update_completed__ps
      -- 
    access_T_CP_0_elements(47) <= access_T_CP_0_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_85_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(46), ack => access_T_CP_0_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	24 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	27 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	26 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_86_sample_start_
      -- 
    access_T_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27);
      gj_access_T_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	24 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	54 
    -- CP-element group 50: 	259 
    -- CP-element group 50: 	265 
    -- CP-element group 50: 	273 
    -- CP-element group 50: 	280 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	28 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_86_update_start_
      -- 
    access_T_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(54) & access_T_CP_0_elements(259) & access_T_CP_0_elements(265) & access_T_CP_0_elements(273) & access_T_CP_0_elements(280);
      gj_access_T_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	26 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_86_sample_start__ps
      -- 
    access_T_CP_0_elements(51) <= access_T_CP_0_elements(26);
    -- CP-element group 52:  join  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	27 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_86_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(52) is bound as output of CP function.
    -- CP-element group 53:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	28 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_86_update_start__ps
      -- 
    access_T_CP_0_elements(53) <= access_T_CP_0_elements(28);
    -- CP-element group 54:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	29 
    -- CP-element group 54: 	259 
    -- CP-element group 54: 	263 
    -- CP-element group 54: 	271 
    -- CP-element group 54: 	279 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	50 
    -- CP-element group 54:  members (15) 
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_index_computed_1
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_index_scaled_1
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_index_resized_1
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_86_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_86_update_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_final_index_sum_regn_Sample/req
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_final_index_sum_regn_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_index_scale_1/scale_rename_ack
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_index_scale_1/scale_rename_req
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_index_scale_1/$exit
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_index_scale_1/$entry
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_index_resize_1/index_resize_ack
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_index_resize_1/index_resize_req
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_index_resize_1/$exit
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_index_resize_1/$entry
      -- 
    req_971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(54), ack => array_obj_ref_269_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(54) is bound as output of CP function.
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	22 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_86_loopback_trigger
      -- 
    access_T_CP_0_elements(55) <= access_T_CP_0_elements(22);
    -- CP-element group 56:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_86_loopback_sample_req
      -- CP-element group 56: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_86_loopback_sample_req_ps
      -- 
    phi_stmt_86_loopback_sample_req_330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_86_loopback_sample_req_330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(56), ack => phi_stmt_86_req_0); -- 
    -- Element group access_T_CP_0_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	23 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_86_entry_trigger
      -- 
    access_T_CP_0_elements(57) <= access_T_CP_0_elements(23);
    -- CP-element group 58:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_86_entry_sample_req
      -- CP-element group 58: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_86_entry_sample_req_ps
      -- 
    phi_stmt_86_entry_sample_req_333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_86_entry_sample_req_333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(58), ack => phi_stmt_86_req_1); -- 
    -- Element group access_T_CP_0_elements(58) is bound as output of CP function.
    -- CP-element group 59:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (2) 
      -- CP-element group 59: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_86_phi_mux_ack
      -- CP-element group 59: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_86_phi_mux_ack_ps
      -- 
    phi_stmt_86_phi_mux_ack_336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_86_ack_0, ack => access_T_CP_0_elements(59)); -- 
    -- CP-element group 60:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (4) 
      -- CP-element group 60: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address2_88_sample_start__ps
      -- CP-element group 60: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address2_88_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address2_88_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address2_88_Sample/req
      -- 
    req_349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(60), ack => n_address2_248_88_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (4) 
      -- CP-element group 61: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address2_88_update_start__ps
      -- CP-element group 61: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address2_88_update_start_
      -- CP-element group 61: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address2_88_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address2_88_Update/req
      -- 
    req_354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(61), ack => n_address2_248_88_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(61) is bound as output of CP function.
    -- CP-element group 62:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address2_88_sample_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address2_88_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address2_88_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address2_88_Sample/ack
      -- 
    ack_350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_248_88_buf_ack_0, ack => access_T_CP_0_elements(62)); -- 
    -- CP-element group 63:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (4) 
      -- CP-element group 63: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address2_88_update_completed__ps
      -- CP-element group 63: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address2_88_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address2_88_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address2_88_Update/ack
      -- 
    ack_355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_248_88_buf_ack_1, ack => access_T_CP_0_elements(63)); -- 
    -- CP-element group 64:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_90_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_90_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_90_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_90_Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_90_sample_start_
      -- 
    rr_367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(66), ack => type_cast_90_inst_req_0); -- 
    access_T_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(64) & access_T_CP_0_elements(68);
      gj_access_T_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_90_update_start_
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_90_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_90_Update/cr
      -- 
    cr_372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(67), ack => type_cast_90_inst_req_1); -- 
    access_T_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(65) & access_T_CP_0_elements(69);
      gj_access_T_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	66 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_90_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_90_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_90_Sample/ra
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_90_sample_completed__ps
      -- 
    ra_368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_90_inst_ack_0, ack => access_T_CP_0_elements(68)); -- 
    -- CP-element group 69:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	67 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_90_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_90_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_90_Update/ca
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_90_update_completed__ps
      -- 
    ca_373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_90_inst_ack_1, ack => access_T_CP_0_elements(69)); -- 
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	24 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	27 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	26 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_91_sample_start_
      -- 
    access_T_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27);
      gj_access_T_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	24 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	75 
    -- CP-element group 71: 	289 
    -- CP-element group 71: 	295 
    -- CP-element group 71: 	303 
    -- CP-element group 71: 	310 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	28 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_91_update_start_
      -- 
    access_T_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(75) & access_T_CP_0_elements(289) & access_T_CP_0_elements(295) & access_T_CP_0_elements(303) & access_T_CP_0_elements(310);
      gj_access_T_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	26 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_91_sample_start__ps
      -- 
    access_T_CP_0_elements(72) <= access_T_CP_0_elements(26);
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	27 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_91_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(73) is bound as output of CP function.
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	28 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_91_update_start__ps
      -- 
    access_T_CP_0_elements(74) <= access_T_CP_0_elements(28);
    -- CP-element group 75:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	29 
    -- CP-element group 75: 	289 
    -- CP-element group 75: 	293 
    -- CP-element group 75: 	301 
    -- CP-element group 75: 	309 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	71 
    -- CP-element group 75:  members (15) 
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_index_scale_1/scale_rename_ack
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_index_scale_1/scale_rename_req
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_index_scale_1/$exit
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_index_scale_1/$entry
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_index_resize_1/index_resize_ack
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_index_resize_1/index_resize_req
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_index_resize_1/$exit
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_index_resize_1/$entry
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_index_computed_1
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_index_scaled_1
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_index_resized_1
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_91_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_91_update_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_final_index_sum_regn_Sample/req
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_final_index_sum_regn_Sample/$entry
      -- 
    req_1137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(75), ack => array_obj_ref_348_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	22 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_91_loopback_trigger
      -- 
    access_T_CP_0_elements(76) <= access_T_CP_0_elements(22);
    -- CP-element group 77:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_91_loopback_sample_req
      -- CP-element group 77: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_91_loopback_sample_req_ps
      -- 
    phi_stmt_91_loopback_sample_req_384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_91_loopback_sample_req_384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(77), ack => phi_stmt_91_req_0); -- 
    -- Element group access_T_CP_0_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	23 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_91_entry_trigger
      -- 
    access_T_CP_0_elements(78) <= access_T_CP_0_elements(23);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_91_entry_sample_req
      -- CP-element group 79: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_91_entry_sample_req_ps
      -- 
    phi_stmt_91_entry_sample_req_387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_91_entry_sample_req_387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(79), ack => phi_stmt_91_req_1); -- 
    -- Element group access_T_CP_0_elements(79) is bound as output of CP function.
    -- CP-element group 80:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_91_phi_mux_ack
      -- CP-element group 80: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_91_phi_mux_ack_ps
      -- 
    phi_stmt_91_phi_mux_ack_390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_91_ack_0, ack => access_T_CP_0_elements(80)); -- 
    -- CP-element group 81:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address3_93_sample_start__ps
      -- CP-element group 81: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address3_93_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address3_93_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address3_93_Sample/req
      -- 
    req_403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(81), ack => n_address3_322_93_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address3_93_update_start__ps
      -- CP-element group 82: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address3_93_update_start_
      -- CP-element group 82: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address3_93_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address3_93_Update/req
      -- 
    req_408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(82), ack => n_address3_322_93_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(82) is bound as output of CP function.
    -- CP-element group 83:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address3_93_sample_completed__ps
      -- CP-element group 83: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address3_93_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address3_93_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address3_93_Sample/ack
      -- 
    ack_404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address3_322_93_buf_ack_0, ack => access_T_CP_0_elements(83)); -- 
    -- CP-element group 84:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address3_93_update_completed__ps
      -- CP-element group 84: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address3_93_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address3_93_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_address3_93_Update/ack
      -- 
    ack_409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address3_322_93_buf_ack_1, ack => access_T_CP_0_elements(84)); -- 
    -- CP-element group 85:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_95_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_95_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: marked-predecessors 
    -- CP-element group 87: 	89 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_95_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_95_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_95_Sample/rr
      -- 
    rr_421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(87), ack => type_cast_95_inst_req_0); -- 
    access_T_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(85) & access_T_CP_0_elements(89);
      gj_access_T_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	90 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_95_update_start_
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_95_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_95_Update/cr
      -- 
    cr_426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(88), ack => type_cast_95_inst_req_1); -- 
    access_T_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(86) & access_T_CP_0_elements(90);
      gj_access_T_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	87 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_95_sample_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_95_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_95_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_95_Sample/ra
      -- 
    ra_422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_0, ack => access_T_CP_0_elements(89)); -- 
    -- CP-element group 90:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	88 
    -- CP-element group 90:  members (4) 
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_95_update_completed__ps
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_95_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_95_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_95_Update/ca
      -- 
    ca_427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_1, ack => access_T_CP_0_elements(90)); -- 
    -- CP-element group 91:  join  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	24 
    -- CP-element group 91: marked-predecessors 
    -- CP-element group 91: 	27 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	26 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_96_sample_start_
      -- 
    access_T_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27);
      gj_access_T_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	24 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	94 
    -- CP-element group 92: 	224 
    -- CP-element group 92: 	254 
    -- CP-element group 92: 	284 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	28 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_96_update_start_
      -- 
    access_T_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(94) & access_T_CP_0_elements(224) & access_T_CP_0_elements(254) & access_T_CP_0_elements(284);
      gj_access_T_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  join  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	27 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_96_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(93) is bound as output of CP function.
    -- CP-element group 94:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	25 
    -- CP-element group 94: 	29 
    -- CP-element group 94: 	222 
    -- CP-element group 94: 	252 
    -- CP-element group 94: 	282 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_96_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_96_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(94) is bound as output of CP function.
    -- CP-element group 95:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	22 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_96_loopback_trigger
      -- 
    access_T_CP_0_elements(95) <= access_T_CP_0_elements(22);
    -- CP-element group 96:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_96_loopback_sample_req
      -- CP-element group 96: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_96_loopback_sample_req_ps
      -- 
    phi_stmt_96_loopback_sample_req_438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_96_loopback_sample_req_438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(96), ack => phi_stmt_96_req_0); -- 
    -- Element group access_T_CP_0_elements(96) is bound as output of CP function.
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	23 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_96_entry_trigger
      -- 
    access_T_CP_0_elements(97) <= access_T_CP_0_elements(23);
    -- CP-element group 98:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_96_entry_sample_req
      -- CP-element group 98: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_96_entry_sample_req_ps
      -- 
    phi_stmt_96_entry_sample_req_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_96_entry_sample_req_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(98), ack => phi_stmt_96_req_1); -- 
    -- Element group access_T_CP_0_elements(98) is bound as output of CP function.
    -- CP-element group 99:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_96_phi_mux_ack
      -- CP-element group 99: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_96_phi_mux_ack_ps
      -- 
    phi_stmt_96_phi_mux_ack_444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_96_ack_0, ack => access_T_CP_0_elements(99)); -- 
    -- CP-element group 100:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (4) 
      -- CP-element group 100: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_mycounter_98_sample_start__ps
      -- CP-element group 100: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_mycounter_98_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_mycounter_98_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_mycounter_98_Sample/req
      -- 
    req_457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(100), ack => n_mycounter_141_98_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_mycounter_98_update_start__ps
      -- CP-element group 101: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_mycounter_98_update_start_
      -- CP-element group 101: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_mycounter_98_Update/$entry
      -- CP-element group 101: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_mycounter_98_Update/req
      -- 
    req_462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(101), ack => n_mycounter_141_98_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(101) is bound as output of CP function.
    -- CP-element group 102:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (4) 
      -- CP-element group 102: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_mycounter_98_sample_completed__ps
      -- CP-element group 102: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_mycounter_98_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_mycounter_98_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_mycounter_98_Sample/ack
      -- 
    ack_458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter_141_98_buf_ack_0, ack => access_T_CP_0_elements(102)); -- 
    -- CP-element group 103:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (4) 
      -- CP-element group 103: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_mycounter_98_update_completed__ps
      -- CP-element group 103: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_mycounter_98_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_mycounter_98_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_mycounter_98_Update/ack
      -- 
    ack_463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter_141_98_buf_ack_1, ack => access_T_CP_0_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (4) 
      -- CP-element group 104: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_100_sample_start__ps
      -- CP-element group 104: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_100_sample_completed__ps
      -- CP-element group 104: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_100_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_100_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(104) is bound as output of CP function.
    -- CP-element group 105:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_100_update_start__ps
      -- CP-element group 105: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_100_update_start_
      -- 
    -- Element group access_T_CP_0_elements(105) is bound as output of CP function.
    -- CP-element group 106:  join  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	107 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_100_update_completed__ps
      -- 
    access_T_CP_0_elements(106) <= access_T_CP_0_elements(107);
    -- CP-element group 107:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	106 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_100_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(107) is a control-delay.
    cp_element_107_delay: control_delay_element  generic map(name => " 107_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(105), ack => access_T_CP_0_elements(107), clk => clk, reset =>reset);
    -- CP-element group 108:  join  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	24 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	27 
    -- CP-element group 108: 	240 
    -- CP-element group 108: 	244 
    -- CP-element group 108: 	248 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	26 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_101_sample_start_
      -- 
    access_T_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27) & access_T_CP_0_elements(240) & access_T_CP_0_elements(244) & access_T_CP_0_elements(248);
      gj_access_T_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	24 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	113 
    -- CP-element group 109: 	247 
    -- CP-element group 109: 	250 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	28 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_101_update_start_
      -- 
    access_T_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(113) & access_T_CP_0_elements(247) & access_T_CP_0_elements(250);
      gj_access_T_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	26 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_101_sample_start__ps
      -- 
    access_T_CP_0_elements(110) <= access_T_CP_0_elements(26);
    -- CP-element group 111:  join  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	27 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_101_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(111) is bound as output of CP function.
    -- CP-element group 112:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	28 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_101_update_start__ps
      -- 
    access_T_CP_0_elements(112) <= access_T_CP_0_elements(28);
    -- CP-element group 113:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	29 
    -- CP-element group 113: 	245 
    -- CP-element group 113: 	249 
    -- CP-element group 113: marked-successors 
    -- CP-element group 113: 	109 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_101_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_101_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(113) is bound as output of CP function.
    -- CP-element group 114:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	22 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_101_loopback_trigger
      -- 
    access_T_CP_0_elements(114) <= access_T_CP_0_elements(22);
    -- CP-element group 115:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_101_loopback_sample_req
      -- CP-element group 115: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_101_loopback_sample_req_ps
      -- 
    phi_stmt_101_loopback_sample_req_482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_101_loopback_sample_req_482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(115), ack => phi_stmt_101_req_0); -- 
    -- Element group access_T_CP_0_elements(115) is bound as output of CP function.
    -- CP-element group 116:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	23 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_101_entry_trigger
      -- 
    access_T_CP_0_elements(116) <= access_T_CP_0_elements(23);
    -- CP-element group 117:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_101_entry_sample_req
      -- CP-element group 117: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_101_entry_sample_req_ps
      -- 
    phi_stmt_101_entry_sample_req_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_101_entry_sample_req_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(117), ack => phi_stmt_101_req_1); -- 
    -- Element group access_T_CP_0_elements(117) is bound as output of CP function.
    -- CP-element group 118:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_101_phi_mux_ack
      -- CP-element group 118: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_101_phi_mux_ack_ps
      -- 
    phi_stmt_101_phi_mux_ack_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_101_ack_0, ack => access_T_CP_0_elements(118)); -- 
    -- CP-element group 119:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (4) 
      -- CP-element group 119: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val1_103_sample_start__ps
      -- CP-element group 119: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val1_103_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val1_103_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val1_103_Sample/req
      -- 
    req_501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(119), ack => n_fetch_val1_217_103_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (4) 
      -- CP-element group 120: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val1_103_update_start__ps
      -- CP-element group 120: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val1_103_update_start_
      -- CP-element group 120: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val1_103_Update/$entry
      -- CP-element group 120: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val1_103_Update/req
      -- 
    req_506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(120), ack => n_fetch_val1_217_103_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(120) is bound as output of CP function.
    -- CP-element group 121:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (4) 
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val1_103_sample_completed__ps
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val1_103_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val1_103_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val1_103_Sample/ack
      -- 
    ack_502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val1_217_103_buf_ack_0, ack => access_T_CP_0_elements(121)); -- 
    -- CP-element group 122:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (4) 
      -- CP-element group 122: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val1_103_update_completed__ps
      -- CP-element group 122: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val1_103_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val1_103_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val1_103_Update/ack
      -- 
    ack_507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val1_217_103_buf_ack_1, ack => access_T_CP_0_elements(122)); -- 
    -- CP-element group 123:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (4) 
      -- CP-element group 123: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch1_104_sample_start__ps
      -- CP-element group 123: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch1_104_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch1_104_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch1_104_Sample/req
      -- 
    req_519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(123), ack => my_fetch1_50_104_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(123) is bound as output of CP function.
    -- CP-element group 124:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (4) 
      -- CP-element group 124: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch1_104_update_start__ps
      -- CP-element group 124: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch1_104_update_start_
      -- CP-element group 124: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch1_104_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch1_104_Update/req
      -- 
    req_524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(124), ack => my_fetch1_50_104_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(124) is bound as output of CP function.
    -- CP-element group 125:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (4) 
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch1_104_sample_completed__ps
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch1_104_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch1_104_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch1_104_Sample/ack
      -- 
    ack_520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch1_50_104_buf_ack_0, ack => access_T_CP_0_elements(125)); -- 
    -- CP-element group 126:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (4) 
      -- CP-element group 126: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch1_104_update_completed__ps
      -- CP-element group 126: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch1_104_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch1_104_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch1_104_Update/ack
      -- 
    ack_525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch1_50_104_buf_ack_1, ack => access_T_CP_0_elements(126)); -- 
    -- CP-element group 127:  join  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	24 
    -- CP-element group 127: marked-predecessors 
    -- CP-element group 127: 	27 
    -- CP-element group 127: 	270 
    -- CP-element group 127: 	274 
    -- CP-element group 127: 	278 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	26 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_105_sample_start_
      -- 
    access_T_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27) & access_T_CP_0_elements(270) & access_T_CP_0_elements(274) & access_T_CP_0_elements(278);
      gj_access_T_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  join  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	24 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	132 
    -- CP-element group 128: 	277 
    -- CP-element group 128: 	280 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	28 
    -- CP-element group 128:  members (1) 
      -- CP-element group 128: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_105_update_start_
      -- 
    access_T_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(132) & access_T_CP_0_elements(277) & access_T_CP_0_elements(280);
      gj_access_T_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	26 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_105_sample_start__ps
      -- 
    access_T_CP_0_elements(129) <= access_T_CP_0_elements(26);
    -- CP-element group 130:  join  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	27 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_105_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(130) is bound as output of CP function.
    -- CP-element group 131:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	28 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_105_update_start__ps
      -- 
    access_T_CP_0_elements(131) <= access_T_CP_0_elements(28);
    -- CP-element group 132:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	29 
    -- CP-element group 132: 	275 
    -- CP-element group 132: 	279 
    -- CP-element group 132: marked-successors 
    -- CP-element group 132: 	128 
    -- CP-element group 132:  members (2) 
      -- CP-element group 132: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_105_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_105_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(132) is bound as output of CP function.
    -- CP-element group 133:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	22 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_105_loopback_trigger
      -- 
    access_T_CP_0_elements(133) <= access_T_CP_0_elements(22);
    -- CP-element group 134:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_105_loopback_sample_req
      -- CP-element group 134: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_105_loopback_sample_req_ps
      -- 
    phi_stmt_105_loopback_sample_req_536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_105_loopback_sample_req_536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(134), ack => phi_stmt_105_req_0); -- 
    -- Element group access_T_CP_0_elements(134) is bound as output of CP function.
    -- CP-element group 135:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	23 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_105_entry_trigger
      -- 
    access_T_CP_0_elements(135) <= access_T_CP_0_elements(23);
    -- CP-element group 136:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (2) 
      -- CP-element group 136: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_105_entry_sample_req
      -- CP-element group 136: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_105_entry_sample_req_ps
      -- 
    phi_stmt_105_entry_sample_req_539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_105_entry_sample_req_539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(136), ack => phi_stmt_105_req_1); -- 
    -- Element group access_T_CP_0_elements(136) is bound as output of CP function.
    -- CP-element group 137:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (2) 
      -- CP-element group 137: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_105_phi_mux_ack
      -- CP-element group 137: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_105_phi_mux_ack_ps
      -- 
    phi_stmt_105_phi_mux_ack_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_105_ack_0, ack => access_T_CP_0_elements(137)); -- 
    -- CP-element group 138:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (4) 
      -- CP-element group 138: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val2_107_sample_start__ps
      -- CP-element group 138: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val2_107_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val2_107_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val2_107_Sample/req
      -- 
    req_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(138), ack => n_fetch_val2_291_107_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(138) is bound as output of CP function.
    -- CP-element group 139:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (4) 
      -- CP-element group 139: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val2_107_update_start__ps
      -- CP-element group 139: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val2_107_update_start_
      -- CP-element group 139: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val2_107_Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val2_107_Update/req
      -- 
    req_560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(139), ack => n_fetch_val2_291_107_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(139) is bound as output of CP function.
    -- CP-element group 140:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val2_107_sample_completed__ps
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val2_107_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val2_107_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val2_107_Sample/ack
      -- 
    ack_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val2_291_107_buf_ack_0, ack => access_T_CP_0_elements(140)); -- 
    -- CP-element group 141:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (4) 
      -- CP-element group 141: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val2_107_update_completed__ps
      -- CP-element group 141: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val2_107_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val2_107_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val2_107_Update/ack
      -- 
    ack_561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val2_291_107_buf_ack_1, ack => access_T_CP_0_elements(141)); -- 
    -- CP-element group 142:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (4) 
      -- CP-element group 142: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch2_108_sample_start__ps
      -- CP-element group 142: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch2_108_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch2_108_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch2_108_Sample/req
      -- 
    req_573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(142), ack => my_fetch2_64_108_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(142) is bound as output of CP function.
    -- CP-element group 143:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (4) 
      -- CP-element group 143: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch2_108_update_start__ps
      -- CP-element group 143: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch2_108_update_start_
      -- CP-element group 143: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch2_108_Update/$entry
      -- CP-element group 143: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch2_108_Update/req
      -- 
    req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(143), ack => my_fetch2_64_108_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(143) is bound as output of CP function.
    -- CP-element group 144:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (4) 
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch2_108_sample_completed__ps
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch2_108_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch2_108_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch2_108_Sample/ack
      -- 
    ack_574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch2_64_108_buf_ack_0, ack => access_T_CP_0_elements(144)); -- 
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (4) 
      -- CP-element group 145: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch2_108_update_completed__ps
      -- CP-element group 145: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch2_108_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch2_108_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch2_108_Update/ack
      -- 
    ack_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch2_64_108_buf_ack_1, ack => access_T_CP_0_elements(145)); -- 
    -- CP-element group 146:  join  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	24 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	27 
    -- CP-element group 146: 	300 
    -- CP-element group 146: 	304 
    -- CP-element group 146: 	308 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	26 
    -- CP-element group 146:  members (1) 
      -- CP-element group 146: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_109_sample_start_
      -- 
    access_T_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27) & access_T_CP_0_elements(300) & access_T_CP_0_elements(304) & access_T_CP_0_elements(308);
      gj_access_T_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  join  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	24 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	151 
    -- CP-element group 147: 	307 
    -- CP-element group 147: 	310 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	28 
    -- CP-element group 147:  members (1) 
      -- CP-element group 147: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_109_update_start_
      -- 
    access_T_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(151) & access_T_CP_0_elements(307) & access_T_CP_0_elements(310);
      gj_access_T_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	26 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_109_sample_start__ps
      -- 
    access_T_CP_0_elements(148) <= access_T_CP_0_elements(26);
    -- CP-element group 149:  join  transition  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	27 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_109_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(149) is bound as output of CP function.
    -- CP-element group 150:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	28 
    -- CP-element group 150: successors 
    -- CP-element group 150:  members (1) 
      -- CP-element group 150: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_109_update_start__ps
      -- 
    access_T_CP_0_elements(150) <= access_T_CP_0_elements(28);
    -- CP-element group 151:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	29 
    -- CP-element group 151: 	305 
    -- CP-element group 151: 	309 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	147 
    -- CP-element group 151:  members (2) 
      -- CP-element group 151: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_109_update_completed_
      -- CP-element group 151: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_109_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(151) is bound as output of CP function.
    -- CP-element group 152:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	22 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (1) 
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_109_loopback_trigger
      -- 
    access_T_CP_0_elements(152) <= access_T_CP_0_elements(22);
    -- CP-element group 153:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (2) 
      -- CP-element group 153: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_109_loopback_sample_req
      -- CP-element group 153: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_109_loopback_sample_req_ps
      -- 
    phi_stmt_109_loopback_sample_req_590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_109_loopback_sample_req_590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(153), ack => phi_stmt_109_req_0); -- 
    -- Element group access_T_CP_0_elements(153) is bound as output of CP function.
    -- CP-element group 154:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	23 
    -- CP-element group 154: successors 
    -- CP-element group 154:  members (1) 
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_109_entry_trigger
      -- 
    access_T_CP_0_elements(154) <= access_T_CP_0_elements(23);
    -- CP-element group 155:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: successors 
    -- CP-element group 155:  members (2) 
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_109_entry_sample_req
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_109_entry_sample_req_ps
      -- 
    phi_stmt_109_entry_sample_req_593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_109_entry_sample_req_593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(155), ack => phi_stmt_109_req_1); -- 
    -- Element group access_T_CP_0_elements(155) is bound as output of CP function.
    -- CP-element group 156:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (2) 
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_109_phi_mux_ack
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_109_phi_mux_ack_ps
      -- 
    phi_stmt_109_phi_mux_ack_596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_109_ack_0, ack => access_T_CP_0_elements(156)); -- 
    -- CP-element group 157:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (4) 
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val3_111_sample_start__ps
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val3_111_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val3_111_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val3_111_Sample/req
      -- 
    req_609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(157), ack => n_fetch_val3_370_111_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(157) is bound as output of CP function.
    -- CP-element group 158:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158:  members (4) 
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val3_111_update_start__ps
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val3_111_update_start_
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val3_111_Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val3_111_Update/req
      -- 
    req_614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(158), ack => n_fetch_val3_370_111_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(158) is bound as output of CP function.
    -- CP-element group 159:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159:  members (4) 
      -- CP-element group 159: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val3_111_sample_completed__ps
      -- CP-element group 159: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val3_111_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val3_111_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val3_111_Sample/ack
      -- 
    ack_610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val3_370_111_buf_ack_0, ack => access_T_CP_0_elements(159)); -- 
    -- CP-element group 160:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (4) 
      -- CP-element group 160: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val3_111_update_completed__ps
      -- CP-element group 160: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val3_111_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val3_111_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_fetch_val3_111_Update/ack
      -- 
    ack_615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_fetch_val3_370_111_buf_ack_1, ack => access_T_CP_0_elements(160)); -- 
    -- CP-element group 161:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (4) 
      -- CP-element group 161: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch3_112_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch3_112_sample_start__ps
      -- CP-element group 161: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch3_112_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch3_112_Sample/req
      -- 
    req_627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(161), ack => my_fetch3_78_112_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(161) is bound as output of CP function.
    -- CP-element group 162:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162:  members (4) 
      -- CP-element group 162: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch3_112_update_start__ps
      -- CP-element group 162: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch3_112_update_start_
      -- CP-element group 162: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch3_112_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch3_112_Update/req
      -- 
    req_632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(162), ack => my_fetch3_78_112_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(162) is bound as output of CP function.
    -- CP-element group 163:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (4) 
      -- CP-element group 163: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch3_112_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch3_112_sample_completed__ps
      -- CP-element group 163: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch3_112_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch3_112_Sample/ack
      -- 
    ack_628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch3_78_112_buf_ack_0, ack => access_T_CP_0_elements(163)); -- 
    -- CP-element group 164:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (4) 
      -- CP-element group 164: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch3_112_update_completed__ps
      -- CP-element group 164: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch3_112_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch3_112_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_my_fetch3_112_Update/ack
      -- 
    ack_633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch3_78_112_buf_ack_1, ack => access_T_CP_0_elements(164)); -- 
    -- CP-element group 165:  join  transition  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	24 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	27 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	26 
    -- CP-element group 165:  members (1) 
      -- CP-element group 165: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_113_sample_start_
      -- 
    access_T_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27);
      gj_access_T_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  join  transition  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	24 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	170 
    -- CP-element group 166: 	224 
    -- CP-element group 166: 	254 
    -- CP-element group 166: 	284 
    -- CP-element group 166: 	310 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	28 
    -- CP-element group 166:  members (1) 
      -- CP-element group 166: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_113_update_start_
      -- 
    access_T_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(170) & access_T_CP_0_elements(224) & access_T_CP_0_elements(254) & access_T_CP_0_elements(284) & access_T_CP_0_elements(310);
      gj_access_T_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	26 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (1) 
      -- CP-element group 167: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_113_sample_start__ps
      -- 
    access_T_CP_0_elements(167) <= access_T_CP_0_elements(26);
    -- CP-element group 168:  join  transition  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	27 
    -- CP-element group 168:  members (1) 
      -- CP-element group 168: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_113_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(168) is bound as output of CP function.
    -- CP-element group 169:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	28 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (1) 
      -- CP-element group 169: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_113_update_start__ps
      -- 
    access_T_CP_0_elements(169) <= access_T_CP_0_elements(28);
    -- CP-element group 170:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	25 
    -- CP-element group 170: 	29 
    -- CP-element group 170: 	222 
    -- CP-element group 170: 	252 
    -- CP-element group 170: 	282 
    -- CP-element group 170: 	309 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	166 
    -- CP-element group 170:  members (2) 
      -- CP-element group 170: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_113_update_completed__ps
      -- CP-element group 170: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_113_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(170) is bound as output of CP function.
    -- CP-element group 171:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	22 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (1) 
      -- CP-element group 171: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_113_loopback_trigger
      -- 
    access_T_CP_0_elements(171) <= access_T_CP_0_elements(22);
    -- CP-element group 172:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (2) 
      -- CP-element group 172: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_113_loopback_sample_req
      -- CP-element group 172: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_113_loopback_sample_req_ps
      -- 
    phi_stmt_113_loopback_sample_req_644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_113_loopback_sample_req_644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(172), ack => phi_stmt_113_req_0); -- 
    -- Element group access_T_CP_0_elements(172) is bound as output of CP function.
    -- CP-element group 173:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	23 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (1) 
      -- CP-element group 173: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_113_entry_trigger
      -- 
    access_T_CP_0_elements(173) <= access_T_CP_0_elements(23);
    -- CP-element group 174:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: successors 
    -- CP-element group 174:  members (2) 
      -- CP-element group 174: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_113_entry_sample_req
      -- CP-element group 174: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_113_entry_sample_req_ps
      -- 
    phi_stmt_113_entry_sample_req_647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_113_entry_sample_req_647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(174), ack => phi_stmt_113_req_1); -- 
    -- Element group access_T_CP_0_elements(174) is bound as output of CP function.
    -- CP-element group 175:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (2) 
      -- CP-element group 175: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_113_phi_mux_ack
      -- CP-element group 175: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_113_phi_mux_ack_ps
      -- 
    phi_stmt_113_phi_mux_ack_650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_113_ack_0, ack => access_T_CP_0_elements(175)); -- 
    -- CP-element group 176:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (4) 
      -- CP-element group 176: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row1_115_sample_start__ps
      -- CP-element group 176: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row1_115_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row1_115_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row1_115_Sample/req
      -- 
    req_663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(176), ack => n_row1_169_115_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(176) is bound as output of CP function.
    -- CP-element group 177:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (4) 
      -- CP-element group 177: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row1_115_update_start__ps
      -- CP-element group 177: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row1_115_update_start_
      -- CP-element group 177: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row1_115_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row1_115_Update/req
      -- 
    req_668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(177), ack => n_row1_169_115_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(177) is bound as output of CP function.
    -- CP-element group 178:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178:  members (4) 
      -- CP-element group 178: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row1_115_sample_completed__ps
      -- CP-element group 178: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row1_115_sample_completed_
      -- CP-element group 178: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row1_115_Sample/$exit
      -- CP-element group 178: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row1_115_Sample/ack
      -- 
    ack_664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row1_169_115_buf_ack_0, ack => access_T_CP_0_elements(178)); -- 
    -- CP-element group 179:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (4) 
      -- CP-element group 179: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row1_115_update_completed__ps
      -- CP-element group 179: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row1_115_update_completed_
      -- CP-element group 179: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row1_115_Update/$exit
      -- CP-element group 179: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row1_115_Update/ack
      -- 
    ack_669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row1_169_115_buf_ack_1, ack => access_T_CP_0_elements(179)); -- 
    -- CP-element group 180:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: successors 
    -- CP-element group 180:  members (4) 
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_117_sample_start__ps
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_117_sample_completed__ps
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_117_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_117_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(180) is bound as output of CP function.
    -- CP-element group 181:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181:  members (2) 
      -- CP-element group 181: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_117_update_start__ps
      -- CP-element group 181: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_117_update_start_
      -- 
    -- Element group access_T_CP_0_elements(181) is bound as output of CP function.
    -- CP-element group 182:  join  transition  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	183 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (1) 
      -- CP-element group 182: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_117_update_completed__ps
      -- 
    access_T_CP_0_elements(182) <= access_T_CP_0_elements(183);
    -- CP-element group 183:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	182 
    -- CP-element group 183:  members (1) 
      -- CP-element group 183: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_117_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(183) is a control-delay.
    cp_element_183_delay: control_delay_element  generic map(name => " 183_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(181), ack => access_T_CP_0_elements(183), clk => clk, reset =>reset);
    -- CP-element group 184:  join  transition  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	24 
    -- CP-element group 184: marked-predecessors 
    -- CP-element group 184: 	27 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	26 
    -- CP-element group 184:  members (1) 
      -- CP-element group 184: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_118_sample_start_
      -- 
    access_T_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27);
      gj_access_T_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  join  transition  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	24 
    -- CP-element group 185: marked-predecessors 
    -- CP-element group 185: 	189 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	28 
    -- CP-element group 185:  members (1) 
      -- CP-element group 185: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_118_update_start_
      -- 
    access_T_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(189);
      gj_access_T_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	26 
    -- CP-element group 186: successors 
    -- CP-element group 186:  members (1) 
      -- CP-element group 186: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_118_sample_start__ps
      -- 
    access_T_CP_0_elements(186) <= access_T_CP_0_elements(26);
    -- CP-element group 187:  join  transition  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	27 
    -- CP-element group 187:  members (1) 
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_118_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(187) is bound as output of CP function.
    -- CP-element group 188:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	28 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (1) 
      -- CP-element group 188: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_118_update_start__ps
      -- 
    access_T_CP_0_elements(188) <= access_T_CP_0_elements(28);
    -- CP-element group 189:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	29 
    -- CP-element group 189: marked-successors 
    -- CP-element group 189: 	185 
    -- CP-element group 189:  members (2) 
      -- CP-element group 189: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_118_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_118_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(189) is bound as output of CP function.
    -- CP-element group 190:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	22 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (1) 
      -- CP-element group 190: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_118_loopback_trigger
      -- 
    access_T_CP_0_elements(190) <= access_T_CP_0_elements(22);
    -- CP-element group 191:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (2) 
      -- CP-element group 191: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_118_loopback_sample_req
      -- CP-element group 191: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_118_loopback_sample_req_ps
      -- 
    phi_stmt_118_loopback_sample_req_688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_118_loopback_sample_req_688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(191), ack => phi_stmt_118_req_1); -- 
    -- Element group access_T_CP_0_elements(191) is bound as output of CP function.
    -- CP-element group 192:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	23 
    -- CP-element group 192: successors 
    -- CP-element group 192:  members (1) 
      -- CP-element group 192: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_118_entry_trigger
      -- 
    access_T_CP_0_elements(192) <= access_T_CP_0_elements(23);
    -- CP-element group 193:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (2) 
      -- CP-element group 193: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_118_entry_sample_req
      -- CP-element group 193: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_118_entry_sample_req_ps
      -- 
    phi_stmt_118_entry_sample_req_691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_118_entry_sample_req_691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(193), ack => phi_stmt_118_req_0); -- 
    -- Element group access_T_CP_0_elements(193) is bound as output of CP function.
    -- CP-element group 194:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (2) 
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_118_phi_mux_ack
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_118_phi_mux_ack_ps
      -- 
    phi_stmt_118_phi_mux_ack_694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_118_ack_0, ack => access_T_CP_0_elements(194)); -- 
    -- CP-element group 195:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (4) 
      -- CP-element group 195: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_121_sample_start__ps
      -- CP-element group 195: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_121_sample_completed__ps
      -- CP-element group 195: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_121_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_121_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(195) is bound as output of CP function.
    -- CP-element group 196:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (2) 
      -- CP-element group 196: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_121_update_start__ps
      -- CP-element group 196: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_121_update_start_
      -- 
    -- Element group access_T_CP_0_elements(196) is bound as output of CP function.
    -- CP-element group 197:  join  transition  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	198 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (1) 
      -- CP-element group 197: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_121_update_completed__ps
      -- 
    access_T_CP_0_elements(197) <= access_T_CP_0_elements(198);
    -- CP-element group 198:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	197 
    -- CP-element group 198:  members (1) 
      -- CP-element group 198: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_121_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(198) is a control-delay.
    cp_element_198_delay: control_delay_element  generic map(name => " 198_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(196), ack => access_T_CP_0_elements(198), clk => clk, reset =>reset);
    -- CP-element group 199:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (4) 
      -- CP-element group 199: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row2_122_sample_start__ps
      -- CP-element group 199: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row2_122_sample_start_
      -- CP-element group 199: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row2_122_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row2_122_Sample/req
      -- 
    req_715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(199), ack => n_row2_243_122_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(199) is bound as output of CP function.
    -- CP-element group 200:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	202 
    -- CP-element group 200:  members (4) 
      -- CP-element group 200: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row2_122_update_start__ps
      -- CP-element group 200: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row2_122_update_start_
      -- CP-element group 200: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row2_122_Update/$entry
      -- CP-element group 200: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row2_122_Update/req
      -- 
    req_720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(200), ack => n_row2_243_122_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(200) is bound as output of CP function.
    -- CP-element group 201:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (4) 
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row2_122_sample_completed__ps
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row2_122_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row2_122_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row2_122_Sample/ack
      -- 
    ack_716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row2_243_122_buf_ack_0, ack => access_T_CP_0_elements(201)); -- 
    -- CP-element group 202:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	200 
    -- CP-element group 202: successors 
    -- CP-element group 202:  members (4) 
      -- CP-element group 202: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row2_122_update_completed__ps
      -- CP-element group 202: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row2_122_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row2_122_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row2_122_Update/ack
      -- 
    ack_721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row2_243_122_buf_ack_1, ack => access_T_CP_0_elements(202)); -- 
    -- CP-element group 203:  join  transition  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	24 
    -- CP-element group 203: marked-predecessors 
    -- CP-element group 203: 	27 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	26 
    -- CP-element group 203:  members (1) 
      -- CP-element group 203: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_123_sample_start_
      -- 
    access_T_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(27);
      gj_access_T_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  join  transition  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	24 
    -- CP-element group 204: marked-predecessors 
    -- CP-element group 204: 	208 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	28 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_123_update_start_
      -- 
    access_T_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(208);
      gj_access_T_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	26 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (1) 
      -- CP-element group 205: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_123_sample_start__ps
      -- 
    access_T_CP_0_elements(205) <= access_T_CP_0_elements(26);
    -- CP-element group 206:  join  transition  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	27 
    -- CP-element group 206:  members (1) 
      -- CP-element group 206: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_123_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(206) is bound as output of CP function.
    -- CP-element group 207:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	28 
    -- CP-element group 207: successors 
    -- CP-element group 207:  members (1) 
      -- CP-element group 207: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_123_update_start__ps
      -- 
    access_T_CP_0_elements(207) <= access_T_CP_0_elements(28);
    -- CP-element group 208:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	29 
    -- CP-element group 208: marked-successors 
    -- CP-element group 208: 	204 
    -- CP-element group 208:  members (2) 
      -- CP-element group 208: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_123_update_completed_
      -- CP-element group 208: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_123_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(208) is bound as output of CP function.
    -- CP-element group 209:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	22 
    -- CP-element group 209: successors 
    -- CP-element group 209:  members (1) 
      -- CP-element group 209: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_123_loopback_trigger
      -- 
    access_T_CP_0_elements(209) <= access_T_CP_0_elements(22);
    -- CP-element group 210:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: successors 
    -- CP-element group 210:  members (2) 
      -- CP-element group 210: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_123_loopback_sample_req
      -- CP-element group 210: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_123_loopback_sample_req_ps
      -- 
    phi_stmt_123_loopback_sample_req_732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_123_loopback_sample_req_732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(210), ack => phi_stmt_123_req_1); -- 
    -- Element group access_T_CP_0_elements(210) is bound as output of CP function.
    -- CP-element group 211:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	23 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (1) 
      -- CP-element group 211: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_123_entry_trigger
      -- 
    access_T_CP_0_elements(211) <= access_T_CP_0_elements(23);
    -- CP-element group 212:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: successors 
    -- CP-element group 212:  members (2) 
      -- CP-element group 212: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_123_entry_sample_req
      -- CP-element group 212: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_123_entry_sample_req_ps
      -- 
    phi_stmt_123_entry_sample_req_735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_123_entry_sample_req_735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(212), ack => phi_stmt_123_req_0); -- 
    -- Element group access_T_CP_0_elements(212) is bound as output of CP function.
    -- CP-element group 213:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (2) 
      -- CP-element group 213: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_123_phi_mux_ack
      -- CP-element group 213: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/phi_stmt_123_phi_mux_ack_ps
      -- 
    phi_stmt_123_phi_mux_ack_738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_123_ack_0, ack => access_T_CP_0_elements(213)); -- 
    -- CP-element group 214:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: successors 
    -- CP-element group 214:  members (4) 
      -- CP-element group 214: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_126_sample_start__ps
      -- CP-element group 214: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_126_sample_completed__ps
      -- CP-element group 214: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_126_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_126_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(214) is bound as output of CP function.
    -- CP-element group 215:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	217 
    -- CP-element group 215:  members (2) 
      -- CP-element group 215: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_126_update_start__ps
      -- CP-element group 215: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_126_update_start_
      -- 
    -- Element group access_T_CP_0_elements(215) is bound as output of CP function.
    -- CP-element group 216:  join  transition  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	217 
    -- CP-element group 216: successors 
    -- CP-element group 216:  members (1) 
      -- CP-element group 216: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_126_update_completed__ps
      -- 
    access_T_CP_0_elements(216) <= access_T_CP_0_elements(217);
    -- CP-element group 217:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	215 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	216 
    -- CP-element group 217:  members (1) 
      -- CP-element group 217: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/type_cast_126_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(217) is a control-delay.
    cp_element_217_delay: control_delay_element  generic map(name => " 217_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(215), ack => access_T_CP_0_elements(217), clk => clk, reset =>reset);
    -- CP-element group 218:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218:  members (4) 
      -- CP-element group 218: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row3_127_sample_start__ps
      -- CP-element group 218: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row3_127_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row3_127_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row3_127_Sample/req
      -- 
    req_759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(218), ack => n_row3_317_127_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(218) is bound as output of CP function.
    -- CP-element group 219:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (4) 
      -- CP-element group 219: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row3_127_update_start__ps
      -- CP-element group 219: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row3_127_update_start_
      -- CP-element group 219: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row3_127_Update/$entry
      -- CP-element group 219: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row3_127_Update/req
      -- 
    req_764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(219), ack => n_row3_317_127_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(219) is bound as output of CP function.
    -- CP-element group 220:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (4) 
      -- CP-element group 220: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row3_127_sample_completed__ps
      -- CP-element group 220: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row3_127_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row3_127_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row3_127_Sample/ack
      -- 
    ack_760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row3_317_127_buf_ack_0, ack => access_T_CP_0_elements(220)); -- 
    -- CP-element group 221:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (4) 
      -- CP-element group 221: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row3_127_update_completed__ps
      -- CP-element group 221: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row3_127_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row3_127_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/R_n_row3_127_Update/ack
      -- 
    ack_765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row3_317_127_buf_ack_1, ack => access_T_CP_0_elements(221)); -- 
    -- CP-element group 222:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	94 
    -- CP-element group 222: 	170 
    -- CP-element group 222: marked-predecessors 
    -- CP-element group 222: 	224 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	224 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_177_sample_start_
      -- CP-element group 222: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_177_Sample/$entry
      -- CP-element group 222: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_177_Sample/req
      -- 
    req_774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(222), ack => W_continue_183_delayed_1_0_175_inst_req_0); -- 
    access_T_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(94) & access_T_CP_0_elements(170) & access_T_CP_0_elements(224);
      gj_access_T_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: marked-predecessors 
    -- CP-element group 223: 	225 
    -- CP-element group 223: 	235 
    -- CP-element group 223: 	243 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_177_update_start_
      -- CP-element group 223: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_177_Update/$entry
      -- CP-element group 223: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_177_Update/req
      -- 
    req_779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(223), ack => W_continue_183_delayed_1_0_175_inst_req_1); -- 
    access_T_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(225) & access_T_CP_0_elements(235) & access_T_CP_0_elements(243);
      gj_access_T_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: successors 
    -- CP-element group 224: marked-successors 
    -- CP-element group 224: 	92 
    -- CP-element group 224: 	166 
    -- CP-element group 224: 	222 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_177_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_177_Sample/$exit
      -- CP-element group 224: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_177_Sample/ack
      -- 
    ack_775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_continue_183_delayed_1_0_175_inst_ack_0, ack => access_T_CP_0_elements(224)); -- 
    -- CP-element group 225:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	233 
    -- CP-element group 225: 	241 
    -- CP-element group 225: marked-successors 
    -- CP-element group 225: 	223 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_177_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_177_Update/$exit
      -- CP-element group 225: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_177_Update/ack
      -- 
    ack_780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_continue_183_delayed_1_0_175_inst_ack_1, ack => access_T_CP_0_elements(225)); -- 
    -- CP-element group 226:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	230 
    -- CP-element group 226: marked-predecessors 
    -- CP-element group 226: 	231 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	231 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_196_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_196_request/$entry
      -- CP-element group 226: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_196_request/req
      -- 
    req_820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(226), ack => addr_of_196_final_reg_req_0); -- 
    access_T_cp_element_group_226: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_226"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(230) & access_T_CP_0_elements(231);
      gj_access_T_cp_element_group_226 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 227:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	24 
    -- CP-element group 227: marked-predecessors 
    -- CP-element group 227: 	232 
    -- CP-element group 227: 	239 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	232 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_196_update_start_
      -- CP-element group 227: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_196_complete/$entry
      -- CP-element group 227: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_196_complete/req
      -- 
    req_825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(227), ack => addr_of_196_final_reg_req_1); -- 
    access_T_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(232) & access_T_CP_0_elements(239);
      gj_access_T_cp_element_group_227 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	24 
    -- CP-element group 228: marked-predecessors 
    -- CP-element group 228: 	230 
    -- CP-element group 228: 	231 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_final_index_sum_regn_update_start
      -- CP-element group 228: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_final_index_sum_regn_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_final_index_sum_regn_Update/req
      -- 
    req_810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(228), ack => array_obj_ref_195_index_offset_req_1); -- 
    access_T_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(230) & access_T_CP_0_elements(231);
      gj_access_T_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	35 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	313 
    -- CP-element group 229: marked-successors 
    -- CP-element group 229: 	31 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_final_index_sum_regn_sample_complete
      -- CP-element group 229: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_final_index_sum_regn_Sample/$exit
      -- CP-element group 229: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_final_index_sum_regn_Sample/ack
      -- 
    ack_806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_195_index_offset_ack_0, ack => access_T_CP_0_elements(229)); -- 
    -- CP-element group 230:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	226 
    -- CP-element group 230: marked-successors 
    -- CP-element group 230: 	228 
    -- CP-element group 230:  members (8) 
      -- CP-element group 230: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_root_address_calculated
      -- CP-element group 230: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_offset_calculated
      -- CP-element group 230: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_final_index_sum_regn_Update/$exit
      -- CP-element group 230: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_final_index_sum_regn_Update/ack
      -- CP-element group 230: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_base_plus_offset/$entry
      -- CP-element group 230: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_base_plus_offset/$exit
      -- CP-element group 230: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_base_plus_offset/sum_rename_req
      -- CP-element group 230: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_195_base_plus_offset/sum_rename_ack
      -- 
    ack_811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_195_index_offset_ack_1, ack => access_T_CP_0_elements(230)); -- 
    -- CP-element group 231:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	226 
    -- CP-element group 231: successors 
    -- CP-element group 231: marked-successors 
    -- CP-element group 231: 	226 
    -- CP-element group 231: 	228 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_196_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_196_request/$exit
      -- CP-element group 231: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_196_request/ack
      -- 
    ack_821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_196_final_reg_ack_0, ack => access_T_CP_0_elements(231)); -- 
    -- CP-element group 232:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	227 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	237 
    -- CP-element group 232: marked-successors 
    -- CP-element group 232: 	227 
    -- CP-element group 232:  members (19) 
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_196_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_196_complete/$exit
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_196_complete/ack
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_base_address_calculated
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_word_address_calculated
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_root_address_calculated
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_base_address_resized
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_base_addr_resize/$entry
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_base_addr_resize/$exit
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_base_addr_resize/base_resize_req
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_base_addr_resize/base_resize_ack
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_base_plus_offset/$entry
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_base_plus_offset/$exit
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_base_plus_offset/sum_rename_req
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_base_plus_offset/sum_rename_ack
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_word_addrgen/$entry
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_word_addrgen/$exit
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_word_addrgen/root_register_req
      -- CP-element group 232: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_word_addrgen/root_register_ack
      -- 
    ack_826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_196_final_reg_ack_1, ack => access_T_CP_0_elements(232)); -- 
    -- CP-element group 233:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	35 
    -- CP-element group 233: 	225 
    -- CP-element group 233: marked-predecessors 
    -- CP-element group 233: 	235 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_200_sample_start_
      -- CP-element group 233: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_200_Sample/$entry
      -- CP-element group 233: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_200_Sample/req
      -- 
    req_834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(233), ack => W_fn1_195_delayed_7_0_198_inst_req_0); -- 
    access_T_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(35) & access_T_CP_0_elements(225) & access_T_CP_0_elements(235);
      gj_access_T_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: marked-predecessors 
    -- CP-element group 234: 	236 
    -- CP-element group 234: 	239 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_200_update_start_
      -- CP-element group 234: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_200_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_200_Update/req
      -- 
    req_839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(234), ack => W_fn1_195_delayed_7_0_198_inst_req_1); -- 
    access_T_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(236) & access_T_CP_0_elements(239);
      gj_access_T_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: marked-successors 
    -- CP-element group 235: 	31 
    -- CP-element group 235: 	223 
    -- CP-element group 235: 	233 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_200_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_200_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_200_Sample/ack
      -- 
    ack_835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn1_195_delayed_7_0_198_inst_ack_0, ack => access_T_CP_0_elements(235)); -- 
    -- CP-element group 236:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236: marked-successors 
    -- CP-element group 236: 	234 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_200_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_200_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_200_Update/ack
      -- 
    ack_840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn1_195_delayed_7_0_198_inst_ack_1, ack => access_T_CP_0_elements(236)); -- 
    -- CP-element group 237:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	232 
    -- CP-element group 237: 	236 
    -- CP-element group 237: marked-predecessors 
    -- CP-element group 237: 	239 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	239 
    -- CP-element group 237:  members (5) 
      -- CP-element group 237: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_sample_start_
      -- CP-element group 237: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Sample/$entry
      -- CP-element group 237: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Sample/word_access_start/$entry
      -- CP-element group 237: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Sample/word_access_start/word_0/$entry
      -- CP-element group 237: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Sample/word_access_start/word_0/rr
      -- 
    rr_873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(237), ack => ptr_deref_204_load_0_req_0); -- 
    access_T_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(232) & access_T_CP_0_elements(236) & access_T_CP_0_elements(239);
      gj_access_T_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	27 
    -- CP-element group 238: marked-predecessors 
    -- CP-element group 238: 	240 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	240 
    -- CP-element group 238:  members (5) 
      -- CP-element group 238: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_update_start_
      -- CP-element group 238: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Update/word_access_complete/$entry
      -- CP-element group 238: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Update/word_access_complete/word_0/$entry
      -- CP-element group 238: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Update/word_access_complete/word_0/cr
      -- 
    cr_884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(238), ack => ptr_deref_204_load_0_req_1); -- 
    access_T_cp_element_group_238: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_238"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(240);
      gj_access_T_cp_element_group_238 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(238), clk => clk, reset => reset); --
    end block;
    -- CP-element group 239:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: successors 
    -- CP-element group 239: marked-successors 
    -- CP-element group 239: 	227 
    -- CP-element group 239: 	234 
    -- CP-element group 239: 	237 
    -- CP-element group 239:  members (5) 
      -- CP-element group 239: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Sample/word_access_start/$exit
      -- CP-element group 239: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Sample/word_access_start/word_0/$exit
      -- CP-element group 239: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Sample/word_access_start/word_0/ra
      -- 
    ra_874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_204_load_0_ack_0, ack => access_T_CP_0_elements(239)); -- 
    -- CP-element group 240:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	313 
    -- CP-element group 240: marked-successors 
    -- CP-element group 240: 	108 
    -- CP-element group 240: 	238 
    -- CP-element group 240:  members (9) 
      -- CP-element group 240: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Update/word_access_complete/$exit
      -- CP-element group 240: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Update/word_access_complete/word_0/$exit
      -- CP-element group 240: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Update/word_access_complete/word_0/ca
      -- CP-element group 240: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Update/ptr_deref_204_Merge/$entry
      -- CP-element group 240: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Update/ptr_deref_204_Merge/$exit
      -- CP-element group 240: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Update/ptr_deref_204_Merge/merge_req
      -- CP-element group 240: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_204_Update/ptr_deref_204_Merge/merge_ack
      -- 
    ca_885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_204_load_0_ack_1, ack => access_T_CP_0_elements(240)); -- 
    -- CP-element group 241:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	35 
    -- CP-element group 241: 	225 
    -- CP-element group 241: marked-predecessors 
    -- CP-element group 241: 	243 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_208_sample_start_
      -- CP-element group 241: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_208_Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_208_Sample/req
      -- 
    req_898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(241), ack => W_fn1_201_delayed_13_0_206_inst_req_0); -- 
    access_T_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(35) & access_T_CP_0_elements(225) & access_T_CP_0_elements(243);
      gj_access_T_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	27 
    -- CP-element group 242: marked-predecessors 
    -- CP-element group 242: 	244 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_208_update_start_
      -- CP-element group 242: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_208_Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_208_Update/req
      -- 
    req_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(242), ack => W_fn1_201_delayed_13_0_206_inst_req_1); -- 
    access_T_cp_element_group_242: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_242"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(244);
      gj_access_T_cp_element_group_242 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(242), clk => clk, reset => reset); --
    end block;
    -- CP-element group 243:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: marked-successors 
    -- CP-element group 243: 	31 
    -- CP-element group 243: 	223 
    -- CP-element group 243: 	241 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_208_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_208_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_208_Sample/ack
      -- 
    ack_899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn1_201_delayed_13_0_206_inst_ack_0, ack => access_T_CP_0_elements(243)); -- 
    -- CP-element group 244:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	313 
    -- CP-element group 244: marked-successors 
    -- CP-element group 244: 	108 
    -- CP-element group 244: 	242 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_208_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_208_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_208_Update/ack
      -- 
    ack_904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn1_201_delayed_13_0_206_inst_ack_1, ack => access_T_CP_0_elements(244)); -- 
    -- CP-element group 245:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	113 
    -- CP-element group 245: marked-predecessors 
    -- CP-element group 245: 	247 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_211_sample_start_
      -- CP-element group 245: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_211_Sample/$entry
      -- CP-element group 245: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_211_Sample/req
      -- 
    req_912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(245), ack => W_fetch_val1_203_delayed_13_0_209_inst_req_0); -- 
    access_T_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(113) & access_T_CP_0_elements(247);
      gj_access_T_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	27 
    -- CP-element group 246: marked-predecessors 
    -- CP-element group 246: 	248 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_211_update_start_
      -- CP-element group 246: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_211_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_211_Update/req
      -- 
    req_917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(246), ack => W_fetch_val1_203_delayed_13_0_209_inst_req_1); -- 
    access_T_cp_element_group_246: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_246"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(248);
      gj_access_T_cp_element_group_246 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(246), clk => clk, reset => reset); --
    end block;
    -- CP-element group 247:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247: marked-successors 
    -- CP-element group 247: 	109 
    -- CP-element group 247: 	245 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_211_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_211_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_211_Sample/ack
      -- 
    ack_913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val1_203_delayed_13_0_209_inst_ack_0, ack => access_T_CP_0_elements(247)); -- 
    -- CP-element group 248:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	313 
    -- CP-element group 248: marked-successors 
    -- CP-element group 248: 	108 
    -- CP-element group 248: 	246 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_211_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_211_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_211_Update/ack
      -- 
    ack_918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val1_203_delayed_13_0_209_inst_ack_1, ack => access_T_CP_0_elements(248)); -- 
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	113 
    -- CP-element group 249: 	35 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	251 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe1_218_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe1_218_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe1_218_Sample/req
      -- 
    req_926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(249), ack => WPIPE_input_pipe1_218_inst_req_0); -- 
    access_T_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(113) & access_T_CP_0_elements(35) & access_T_CP_0_elements(251);
      gj_access_T_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250: marked-successors 
    -- CP-element group 250: 	109 
    -- CP-element group 250: 	31 
    -- CP-element group 250:  members (6) 
      -- CP-element group 250: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe1_218_sample_completed_
      -- CP-element group 250: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe1_218_update_start_
      -- CP-element group 250: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe1_218_Sample/$exit
      -- CP-element group 250: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe1_218_Sample/ack
      -- CP-element group 250: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe1_218_Update/$entry
      -- CP-element group 250: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe1_218_Update/req
      -- 
    ack_927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_218_inst_ack_0, ack => access_T_CP_0_elements(250)); -- 
    req_931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(250), ack => WPIPE_input_pipe1_218_inst_req_1); -- 
    -- CP-element group 251:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	313 
    -- CP-element group 251: marked-successors 
    -- CP-element group 251: 	249 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe1_218_update_completed_
      -- CP-element group 251: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe1_218_Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe1_218_Update/ack
      -- 
    ack_932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_218_inst_ack_1, ack => access_T_CP_0_elements(251)); -- 
    -- CP-element group 252:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	94 
    -- CP-element group 252: 	170 
    -- CP-element group 252: marked-predecessors 
    -- CP-element group 252: 	254 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	254 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_251_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_251_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_251_Sample/req
      -- 
    req_940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(252), ack => W_continue_245_delayed_1_0_249_inst_req_0); -- 
    access_T_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(94) & access_T_CP_0_elements(170) & access_T_CP_0_elements(254);
      gj_access_T_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: marked-predecessors 
    -- CP-element group 253: 	255 
    -- CP-element group 253: 	265 
    -- CP-element group 253: 	273 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_251_update_start_
      -- CP-element group 253: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_251_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_251_Update/req
      -- 
    req_945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(253), ack => W_continue_245_delayed_1_0_249_inst_req_1); -- 
    access_T_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(255) & access_T_CP_0_elements(265) & access_T_CP_0_elements(273);
      gj_access_T_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	252 
    -- CP-element group 254: successors 
    -- CP-element group 254: marked-successors 
    -- CP-element group 254: 	92 
    -- CP-element group 254: 	166 
    -- CP-element group 254: 	252 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_251_sample_completed_
      -- CP-element group 254: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_251_Sample/$exit
      -- CP-element group 254: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_251_Sample/ack
      -- 
    ack_941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_continue_245_delayed_1_0_249_inst_ack_0, ack => access_T_CP_0_elements(254)); -- 
    -- CP-element group 255:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	263 
    -- CP-element group 255: 	271 
    -- CP-element group 255: marked-successors 
    -- CP-element group 255: 	253 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_251_update_completed_
      -- CP-element group 255: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_251_Update/$exit
      -- CP-element group 255: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_251_Update/ack
      -- 
    ack_946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_continue_245_delayed_1_0_249_inst_ack_1, ack => access_T_CP_0_elements(255)); -- 
    -- CP-element group 256:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	260 
    -- CP-element group 256: marked-predecessors 
    -- CP-element group 256: 	261 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	261 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_270_request/req
      -- CP-element group 256: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_270_request/$entry
      -- CP-element group 256: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_270_sample_start_
      -- 
    req_986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(256), ack => addr_of_270_final_reg_req_0); -- 
    access_T_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(260) & access_T_CP_0_elements(261);
      gj_access_T_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	24 
    -- CP-element group 257: marked-predecessors 
    -- CP-element group 257: 	262 
    -- CP-element group 257: 	269 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	262 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_270_complete/req
      -- CP-element group 257: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_270_complete/$entry
      -- CP-element group 257: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_270_update_start_
      -- 
    req_991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(257), ack => addr_of_270_final_reg_req_1); -- 
    access_T_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(262) & access_T_CP_0_elements(269);
      gj_access_T_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	24 
    -- CP-element group 258: marked-predecessors 
    -- CP-element group 258: 	260 
    -- CP-element group 258: 	261 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	260 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_final_index_sum_regn_Update/req
      -- CP-element group 258: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_final_index_sum_regn_Update/$entry
      -- CP-element group 258: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_final_index_sum_regn_update_start
      -- 
    req_976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(258), ack => array_obj_ref_269_index_offset_req_1); -- 
    access_T_cp_element_group_258: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_258"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(260) & access_T_CP_0_elements(261);
      gj_access_T_cp_element_group_258 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(258), clk => clk, reset => reset); --
    end block;
    -- CP-element group 259:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	54 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	313 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	50 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_final_index_sum_regn_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_final_index_sum_regn_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_final_index_sum_regn_sample_complete
      -- 
    ack_972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_269_index_offset_ack_0, ack => access_T_CP_0_elements(259)); -- 
    -- CP-element group 260:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	256 
    -- CP-element group 260: marked-successors 
    -- CP-element group 260: 	258 
    -- CP-element group 260:  members (8) 
      -- CP-element group 260: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_offset_calculated
      -- CP-element group 260: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_base_plus_offset/$exit
      -- CP-element group 260: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_base_plus_offset/sum_rename_ack
      -- CP-element group 260: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_base_plus_offset/sum_rename_req
      -- CP-element group 260: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_root_address_calculated
      -- CP-element group 260: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_base_plus_offset/$entry
      -- CP-element group 260: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_final_index_sum_regn_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_269_final_index_sum_regn_Update/$exit
      -- 
    ack_977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_269_index_offset_ack_1, ack => access_T_CP_0_elements(260)); -- 
    -- CP-element group 261:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	256 
    -- CP-element group 261: successors 
    -- CP-element group 261: marked-successors 
    -- CP-element group 261: 	256 
    -- CP-element group 261: 	258 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_270_request/ack
      -- CP-element group 261: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_270_request/$exit
      -- CP-element group 261: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_270_sample_completed_
      -- 
    ack_987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_270_final_reg_ack_0, ack => access_T_CP_0_elements(261)); -- 
    -- CP-element group 262:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	257 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	267 
    -- CP-element group 262: marked-successors 
    -- CP-element group 262: 	257 
    -- CP-element group 262:  members (19) 
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_270_update_completed_
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_270_complete/ack
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_270_complete/$exit
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_word_addrgen/root_register_ack
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_word_addrgen/root_register_req
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_word_addrgen/$exit
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_word_addrgen/$entry
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_base_plus_offset/sum_rename_ack
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_base_plus_offset/sum_rename_req
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_base_plus_offset/$exit
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_base_plus_offset/$entry
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_base_addr_resize/base_resize_ack
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_base_addr_resize/base_resize_req
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_base_addr_resize/$exit
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_base_addr_resize/$entry
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_base_address_resized
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_root_address_calculated
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_word_address_calculated
      -- CP-element group 262: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_base_address_calculated
      -- 
    ack_992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_270_final_reg_ack_1, ack => access_T_CP_0_elements(262)); -- 
    -- CP-element group 263:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	54 
    -- CP-element group 263: 	255 
    -- CP-element group 263: marked-predecessors 
    -- CP-element group 263: 	265 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	265 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_274_Sample/req
      -- CP-element group 263: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_274_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_274_sample_start_
      -- 
    req_1000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(263), ack => W_fn2_257_delayed_7_0_272_inst_req_0); -- 
    access_T_cp_element_group_263: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_263"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(54) & access_T_CP_0_elements(255) & access_T_CP_0_elements(265);
      gj_access_T_cp_element_group_263 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(263), clk => clk, reset => reset); --
    end block;
    -- CP-element group 264:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: marked-predecessors 
    -- CP-element group 264: 	266 
    -- CP-element group 264: 	269 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	266 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_274_Update/req
      -- CP-element group 264: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_274_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_274_update_start_
      -- 
    req_1005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(264), ack => W_fn2_257_delayed_7_0_272_inst_req_1); -- 
    access_T_cp_element_group_264: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_264"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(266) & access_T_CP_0_elements(269);
      gj_access_T_cp_element_group_264 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(264), clk => clk, reset => reset); --
    end block;
    -- CP-element group 265:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	263 
    -- CP-element group 265: successors 
    -- CP-element group 265: marked-successors 
    -- CP-element group 265: 	50 
    -- CP-element group 265: 	253 
    -- CP-element group 265: 	263 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_274_Sample/ack
      -- CP-element group 265: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_274_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_274_sample_completed_
      -- 
    ack_1001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn2_257_delayed_7_0_272_inst_ack_0, ack => access_T_CP_0_elements(265)); -- 
    -- CP-element group 266:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	264 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266: marked-successors 
    -- CP-element group 266: 	264 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_274_Update/ack
      -- CP-element group 266: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_274_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_274_update_completed_
      -- 
    ack_1006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn2_257_delayed_7_0_272_inst_ack_1, ack => access_T_CP_0_elements(266)); -- 
    -- CP-element group 267:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	262 
    -- CP-element group 267: 	266 
    -- CP-element group 267: marked-predecessors 
    -- CP-element group 267: 	269 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	269 
    -- CP-element group 267:  members (5) 
      -- CP-element group 267: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Sample/word_access_start/word_0/rr
      -- CP-element group 267: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Sample/word_access_start/word_0/$entry
      -- CP-element group 267: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Sample/word_access_start/$entry
      -- CP-element group 267: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_sample_start_
      -- 
    rr_1039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(267), ack => ptr_deref_278_load_0_req_0); -- 
    access_T_cp_element_group_267: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_267"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(262) & access_T_CP_0_elements(266) & access_T_CP_0_elements(269);
      gj_access_T_cp_element_group_267 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(267), clk => clk, reset => reset); --
    end block;
    -- CP-element group 268:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	27 
    -- CP-element group 268: marked-predecessors 
    -- CP-element group 268: 	270 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	270 
    -- CP-element group 268:  members (5) 
      -- CP-element group 268: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Update/word_access_complete/word_0/cr
      -- CP-element group 268: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Update/word_access_complete/word_0/$entry
      -- CP-element group 268: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Update/word_access_complete/$entry
      -- CP-element group 268: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Update/$entry
      -- CP-element group 268: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_update_start_
      -- 
    cr_1050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(268), ack => ptr_deref_278_load_0_req_1); -- 
    access_T_cp_element_group_268: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_268"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(270);
      gj_access_T_cp_element_group_268 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(268), clk => clk, reset => reset); --
    end block;
    -- CP-element group 269:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	267 
    -- CP-element group 269: successors 
    -- CP-element group 269: marked-successors 
    -- CP-element group 269: 	257 
    -- CP-element group 269: 	264 
    -- CP-element group 269: 	267 
    -- CP-element group 269:  members (5) 
      -- CP-element group 269: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Sample/word_access_start/word_0/ra
      -- CP-element group 269: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Sample/word_access_start/word_0/$exit
      -- CP-element group 269: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Sample/word_access_start/$exit
      -- CP-element group 269: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_sample_completed_
      -- 
    ra_1040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_278_load_0_ack_0, ack => access_T_CP_0_elements(269)); -- 
    -- CP-element group 270:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	268 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	313 
    -- CP-element group 270: marked-successors 
    -- CP-element group 270: 	127 
    -- CP-element group 270: 	268 
    -- CP-element group 270:  members (9) 
      -- CP-element group 270: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Update/ptr_deref_278_Merge/merge_ack
      -- CP-element group 270: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Update/ptr_deref_278_Merge/merge_req
      -- CP-element group 270: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Update/ptr_deref_278_Merge/$exit
      -- CP-element group 270: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Update/ptr_deref_278_Merge/$entry
      -- CP-element group 270: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Update/word_access_complete/word_0/ca
      -- CP-element group 270: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Update/word_access_complete/word_0/$exit
      -- CP-element group 270: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Update/word_access_complete/$exit
      -- CP-element group 270: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_278_update_completed_
      -- 
    ca_1051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_278_load_0_ack_1, ack => access_T_CP_0_elements(270)); -- 
    -- CP-element group 271:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	54 
    -- CP-element group 271: 	255 
    -- CP-element group 271: marked-predecessors 
    -- CP-element group 271: 	273 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	273 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_282_Sample/req
      -- CP-element group 271: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_282_Sample/$entry
      -- CP-element group 271: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_282_sample_start_
      -- 
    req_1064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(271), ack => W_fn2_263_delayed_13_0_280_inst_req_0); -- 
    access_T_cp_element_group_271: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_271"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(54) & access_T_CP_0_elements(255) & access_T_CP_0_elements(273);
      gj_access_T_cp_element_group_271 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(271), clk => clk, reset => reset); --
    end block;
    -- CP-element group 272:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	27 
    -- CP-element group 272: marked-predecessors 
    -- CP-element group 272: 	274 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	274 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_282_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_282_update_start_
      -- CP-element group 272: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_282_Update/req
      -- 
    req_1069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(272), ack => W_fn2_263_delayed_13_0_280_inst_req_1); -- 
    access_T_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(274);
      gj_access_T_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	271 
    -- CP-element group 273: successors 
    -- CP-element group 273: marked-successors 
    -- CP-element group 273: 	50 
    -- CP-element group 273: 	253 
    -- CP-element group 273: 	271 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_282_Sample/ack
      -- CP-element group 273: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_282_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_282_sample_completed_
      -- 
    ack_1065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn2_263_delayed_13_0_280_inst_ack_0, ack => access_T_CP_0_elements(273)); -- 
    -- CP-element group 274:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	272 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	313 
    -- CP-element group 274: marked-successors 
    -- CP-element group 274: 	127 
    -- CP-element group 274: 	272 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_282_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_282_update_completed_
      -- CP-element group 274: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_282_Update/ack
      -- 
    ack_1070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn2_263_delayed_13_0_280_inst_ack_1, ack => access_T_CP_0_elements(274)); -- 
    -- CP-element group 275:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	132 
    -- CP-element group 275: marked-predecessors 
    -- CP-element group 275: 	277 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	277 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_285_Sample/$entry
      -- CP-element group 275: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_285_sample_start_
      -- CP-element group 275: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_285_Sample/req
      -- 
    req_1078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(275), ack => W_fetch_val2_265_delayed_13_0_283_inst_req_0); -- 
    access_T_cp_element_group_275: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_275"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(132) & access_T_CP_0_elements(277);
      gj_access_T_cp_element_group_275 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(275), clk => clk, reset => reset); --
    end block;
    -- CP-element group 276:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	27 
    -- CP-element group 276: marked-predecessors 
    -- CP-element group 276: 	278 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	278 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_285_update_start_
      -- CP-element group 276: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_285_Update/req
      -- CP-element group 276: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_285_Update/$entry
      -- 
    req_1083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(276), ack => W_fetch_val2_265_delayed_13_0_283_inst_req_1); -- 
    access_T_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(278);
      gj_access_T_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	275 
    -- CP-element group 277: successors 
    -- CP-element group 277: marked-successors 
    -- CP-element group 277: 	128 
    -- CP-element group 277: 	275 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_285_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_285_sample_completed_
      -- CP-element group 277: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_285_Sample/ack
      -- 
    ack_1079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val2_265_delayed_13_0_283_inst_ack_0, ack => access_T_CP_0_elements(277)); -- 
    -- CP-element group 278:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	276 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	313 
    -- CP-element group 278: marked-successors 
    -- CP-element group 278: 	127 
    -- CP-element group 278: 	276 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_285_update_completed_
      -- CP-element group 278: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_285_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_285_Update/$exit
      -- 
    ack_1084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val2_265_delayed_13_0_283_inst_ack_1, ack => access_T_CP_0_elements(278)); -- 
    -- CP-element group 279:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	54 
    -- CP-element group 279: 	132 
    -- CP-element group 279: marked-predecessors 
    -- CP-element group 279: 	281 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe2_292_Sample/req
      -- CP-element group 279: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe2_292_Sample/$entry
      -- CP-element group 279: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe2_292_sample_start_
      -- 
    req_1092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(279), ack => WPIPE_input_pipe2_292_inst_req_0); -- 
    access_T_cp_element_group_279: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_279"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(54) & access_T_CP_0_elements(132) & access_T_CP_0_elements(281);
      gj_access_T_cp_element_group_279 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(279), clk => clk, reset => reset); --
    end block;
    -- CP-element group 280:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280: marked-successors 
    -- CP-element group 280: 	50 
    -- CP-element group 280: 	128 
    -- CP-element group 280:  members (6) 
      -- CP-element group 280: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe2_292_Update/req
      -- CP-element group 280: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe2_292_Update/$entry
      -- CP-element group 280: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe2_292_Sample/ack
      -- CP-element group 280: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe2_292_Sample/$exit
      -- CP-element group 280: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe2_292_update_start_
      -- CP-element group 280: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe2_292_sample_completed_
      -- 
    ack_1093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe2_292_inst_ack_0, ack => access_T_CP_0_elements(280)); -- 
    req_1097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(280), ack => WPIPE_input_pipe2_292_inst_req_1); -- 
    -- CP-element group 281:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	313 
    -- CP-element group 281: marked-successors 
    -- CP-element group 281: 	279 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe2_292_Update/ack
      -- CP-element group 281: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe2_292_Update/$exit
      -- CP-element group 281: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe2_292_update_completed_
      -- 
    ack_1098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe2_292_inst_ack_1, ack => access_T_CP_0_elements(281)); -- 
    -- CP-element group 282:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	94 
    -- CP-element group 282: 	170 
    -- CP-element group 282: marked-predecessors 
    -- CP-element group 282: 	284 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	284 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_325_Sample/req
      -- CP-element group 282: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_325_Sample/$entry
      -- CP-element group 282: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_325_sample_start_
      -- 
    req_1106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(282), ack => W_continue_307_delayed_1_0_323_inst_req_0); -- 
    access_T_cp_element_group_282: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_282"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(94) & access_T_CP_0_elements(170) & access_T_CP_0_elements(284);
      gj_access_T_cp_element_group_282 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(282), clk => clk, reset => reset); --
    end block;
    -- CP-element group 283:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: marked-predecessors 
    -- CP-element group 283: 	285 
    -- CP-element group 283: 	295 
    -- CP-element group 283: 	303 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	285 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_325_Update/req
      -- CP-element group 283: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_325_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_325_update_start_
      -- 
    req_1111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(283), ack => W_continue_307_delayed_1_0_323_inst_req_1); -- 
    access_T_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(285) & access_T_CP_0_elements(295) & access_T_CP_0_elements(303);
      gj_access_T_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	282 
    -- CP-element group 284: successors 
    -- CP-element group 284: marked-successors 
    -- CP-element group 284: 	92 
    -- CP-element group 284: 	166 
    -- CP-element group 284: 	282 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_325_Sample/ack
      -- CP-element group 284: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_325_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_325_sample_completed_
      -- 
    ack_1107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_continue_307_delayed_1_0_323_inst_ack_0, ack => access_T_CP_0_elements(284)); -- 
    -- CP-element group 285:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	283 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	293 
    -- CP-element group 285: 	301 
    -- CP-element group 285: marked-successors 
    -- CP-element group 285: 	283 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_325_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_325_update_completed_
      -- CP-element group 285: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_325_Update/ack
      -- 
    ack_1112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_continue_307_delayed_1_0_323_inst_ack_1, ack => access_T_CP_0_elements(285)); -- 
    -- CP-element group 286:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	290 
    -- CP-element group 286: marked-predecessors 
    -- CP-element group 286: 	291 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	291 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_349_request/req
      -- CP-element group 286: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_349_request/$entry
      -- CP-element group 286: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_349_sample_start_
      -- 
    req_1152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(286), ack => addr_of_349_final_reg_req_0); -- 
    access_T_cp_element_group_286: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_286"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(290) & access_T_CP_0_elements(291);
      gj_access_T_cp_element_group_286 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(286), clk => clk, reset => reset); --
    end block;
    -- CP-element group 287:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	24 
    -- CP-element group 287: marked-predecessors 
    -- CP-element group 287: 	292 
    -- CP-element group 287: 	299 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	292 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_349_complete/$entry
      -- CP-element group 287: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_349_update_start_
      -- CP-element group 287: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_349_complete/req
      -- 
    req_1157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(287), ack => addr_of_349_final_reg_req_1); -- 
    access_T_cp_element_group_287: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_287"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(292) & access_T_CP_0_elements(299);
      gj_access_T_cp_element_group_287 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(287), clk => clk, reset => reset); --
    end block;
    -- CP-element group 288:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	24 
    -- CP-element group 288: marked-predecessors 
    -- CP-element group 288: 	290 
    -- CP-element group 288: 	291 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	290 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_final_index_sum_regn_Update/req
      -- CP-element group 288: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_final_index_sum_regn_Update/$entry
      -- CP-element group 288: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_final_index_sum_regn_update_start
      -- 
    req_1142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(288), ack => array_obj_ref_348_index_offset_req_1); -- 
    access_T_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(24) & access_T_CP_0_elements(290) & access_T_CP_0_elements(291);
      gj_access_T_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	75 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	313 
    -- CP-element group 289: marked-successors 
    -- CP-element group 289: 	71 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_final_index_sum_regn_Sample/ack
      -- CP-element group 289: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_final_index_sum_regn_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_final_index_sum_regn_sample_complete
      -- 
    ack_1138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_348_index_offset_ack_0, ack => access_T_CP_0_elements(289)); -- 
    -- CP-element group 290:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	288 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	286 
    -- CP-element group 290: marked-successors 
    -- CP-element group 290: 	288 
    -- CP-element group 290:  members (8) 
      -- CP-element group 290: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_base_plus_offset/sum_rename_ack
      -- CP-element group 290: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_offset_calculated
      -- CP-element group 290: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_root_address_calculated
      -- CP-element group 290: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_base_plus_offset/sum_rename_req
      -- CP-element group 290: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_base_plus_offset/$exit
      -- CP-element group 290: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_base_plus_offset/$entry
      -- CP-element group 290: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_final_index_sum_regn_Update/ack
      -- CP-element group 290: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/array_obj_ref_348_final_index_sum_regn_Update/$exit
      -- 
    ack_1143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_348_index_offset_ack_1, ack => access_T_CP_0_elements(290)); -- 
    -- CP-element group 291:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	286 
    -- CP-element group 291: successors 
    -- CP-element group 291: marked-successors 
    -- CP-element group 291: 	286 
    -- CP-element group 291: 	288 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_349_request/$exit
      -- CP-element group 291: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_349_request/ack
      -- CP-element group 291: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_349_sample_completed_
      -- 
    ack_1153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_349_final_reg_ack_0, ack => access_T_CP_0_elements(291)); -- 
    -- CP-element group 292:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	287 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	297 
    -- CP-element group 292: marked-successors 
    -- CP-element group 292: 	287 
    -- CP-element group 292:  members (19) 
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_349_complete/$exit
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_root_address_calculated
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_word_addrgen/$entry
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_base_address_resized
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_word_addrgen/root_register_ack
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_word_addrgen/root_register_req
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_word_addrgen/$exit
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_word_address_calculated
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_base_address_calculated
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_base_plus_offset/sum_rename_ack
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_base_plus_offset/sum_rename_req
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_base_plus_offset/$exit
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_349_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_base_plus_offset/$entry
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/addr_of_349_complete/ack
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_base_addr_resize/base_resize_ack
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_base_addr_resize/base_resize_req
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_base_addr_resize/$exit
      -- CP-element group 292: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_base_addr_resize/$entry
      -- 
    ack_1158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_349_final_reg_ack_1, ack => access_T_CP_0_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	75 
    -- CP-element group 293: 	285 
    -- CP-element group 293: marked-predecessors 
    -- CP-element group 293: 	295 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	295 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_353_sample_start_
      -- CP-element group 293: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_353_Sample/req
      -- CP-element group 293: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_353_Sample/$entry
      -- 
    req_1166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(293), ack => W_fn3_324_delayed_7_0_351_inst_req_0); -- 
    access_T_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(75) & access_T_CP_0_elements(285) & access_T_CP_0_elements(295);
      gj_access_T_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: marked-predecessors 
    -- CP-element group 294: 	296 
    -- CP-element group 294: 	299 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	296 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_353_Update/req
      -- CP-element group 294: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_353_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_353_update_start_
      -- 
    req_1171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(294), ack => W_fn3_324_delayed_7_0_351_inst_req_1); -- 
    access_T_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(296) & access_T_CP_0_elements(299);
      gj_access_T_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	293 
    -- CP-element group 295: successors 
    -- CP-element group 295: marked-successors 
    -- CP-element group 295: 	71 
    -- CP-element group 295: 	283 
    -- CP-element group 295: 	293 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_353_sample_completed_
      -- CP-element group 295: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_353_Sample/ack
      -- CP-element group 295: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_353_Sample/$exit
      -- 
    ack_1167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn3_324_delayed_7_0_351_inst_ack_0, ack => access_T_CP_0_elements(295)); -- 
    -- CP-element group 296:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	294 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296: marked-successors 
    -- CP-element group 296: 	294 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_353_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_353_update_completed_
      -- CP-element group 296: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_353_Update/ack
      -- 
    ack_1172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn3_324_delayed_7_0_351_inst_ack_1, ack => access_T_CP_0_elements(296)); -- 
    -- CP-element group 297:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	292 
    -- CP-element group 297: 	296 
    -- CP-element group 297: marked-predecessors 
    -- CP-element group 297: 	299 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	299 
    -- CP-element group 297:  members (5) 
      -- CP-element group 297: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Sample/word_access_start/word_0/$entry
      -- CP-element group 297: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Sample/word_access_start/$entry
      -- CP-element group 297: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Sample/$entry
      -- CP-element group 297: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_sample_start_
      -- CP-element group 297: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Sample/word_access_start/word_0/rr
      -- 
    rr_1205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(297), ack => ptr_deref_357_load_0_req_0); -- 
    access_T_cp_element_group_297: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_297"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(292) & access_T_CP_0_elements(296) & access_T_CP_0_elements(299);
      gj_access_T_cp_element_group_297 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(297), clk => clk, reset => reset); --
    end block;
    -- CP-element group 298:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	27 
    -- CP-element group 298: marked-predecessors 
    -- CP-element group 298: 	300 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	300 
    -- CP-element group 298:  members (5) 
      -- CP-element group 298: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Update/word_access_complete/word_0/cr
      -- CP-element group 298: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Update/word_access_complete/word_0/$entry
      -- CP-element group 298: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Update/word_access_complete/$entry
      -- CP-element group 298: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_update_start_
      -- 
    cr_1216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(298), ack => ptr_deref_357_load_0_req_1); -- 
    access_T_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(300);
      gj_access_T_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	297 
    -- CP-element group 299: successors 
    -- CP-element group 299: marked-successors 
    -- CP-element group 299: 	287 
    -- CP-element group 299: 	294 
    -- CP-element group 299: 	297 
    -- CP-element group 299:  members (5) 
      -- CP-element group 299: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Sample/word_access_start/$exit
      -- CP-element group 299: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Sample/word_access_start/word_0/ra
      -- CP-element group 299: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Sample/word_access_start/word_0/$exit
      -- 
    ra_1206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_357_load_0_ack_0, ack => access_T_CP_0_elements(299)); -- 
    -- CP-element group 300:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	298 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	313 
    -- CP-element group 300: marked-successors 
    -- CP-element group 300: 	146 
    -- CP-element group 300: 	298 
    -- CP-element group 300:  members (9) 
      -- CP-element group 300: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Update/ptr_deref_357_Merge/merge_ack
      -- CP-element group 300: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Update/word_access_complete/word_0/$exit
      -- CP-element group 300: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Update/ptr_deref_357_Merge/merge_req
      -- CP-element group 300: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Update/word_access_complete/$exit
      -- CP-element group 300: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Update/ptr_deref_357_Merge/$entry
      -- CP-element group 300: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Update/ptr_deref_357_Merge/$exit
      -- CP-element group 300: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/ptr_deref_357_Update/word_access_complete/word_0/ca
      -- 
    ca_1217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_357_load_0_ack_1, ack => access_T_CP_0_elements(300)); -- 
    -- CP-element group 301:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	75 
    -- CP-element group 301: 	285 
    -- CP-element group 301: marked-predecessors 
    -- CP-element group 301: 	303 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	303 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_361_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_361_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_361_Sample/req
      -- 
    req_1230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(301), ack => W_fn3_330_delayed_13_0_359_inst_req_0); -- 
    access_T_cp_element_group_301: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_301"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(75) & access_T_CP_0_elements(285) & access_T_CP_0_elements(303);
      gj_access_T_cp_element_group_301 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(301), clk => clk, reset => reset); --
    end block;
    -- CP-element group 302:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	27 
    -- CP-element group 302: marked-predecessors 
    -- CP-element group 302: 	304 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	304 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_361_Update/req
      -- CP-element group 302: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_361_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_361_update_start_
      -- 
    req_1235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(302), ack => W_fn3_330_delayed_13_0_359_inst_req_1); -- 
    access_T_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(304);
      gj_access_T_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	301 
    -- CP-element group 303: successors 
    -- CP-element group 303: marked-successors 
    -- CP-element group 303: 	71 
    -- CP-element group 303: 	283 
    -- CP-element group 303: 	301 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_361_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_361_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_361_sample_completed_
      -- 
    ack_1231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn3_330_delayed_13_0_359_inst_ack_0, ack => access_T_CP_0_elements(303)); -- 
    -- CP-element group 304:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	302 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	313 
    -- CP-element group 304: marked-successors 
    -- CP-element group 304: 	146 
    -- CP-element group 304: 	302 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_361_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_361_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_361_Update/$exit
      -- 
    ack_1236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn3_330_delayed_13_0_359_inst_ack_1, ack => access_T_CP_0_elements(304)); -- 
    -- CP-element group 305:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	151 
    -- CP-element group 305: marked-predecessors 
    -- CP-element group 305: 	307 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_364_Sample/req
      -- CP-element group 305: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_364_sample_start_
      -- CP-element group 305: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_364_Sample/$entry
      -- 
    req_1244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(305), ack => W_fetch_val3_332_delayed_13_0_362_inst_req_0); -- 
    access_T_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(151) & access_T_CP_0_elements(307);
      gj_access_T_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	27 
    -- CP-element group 306: marked-predecessors 
    -- CP-element group 306: 	308 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	308 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_364_Update/req
      -- CP-element group 306: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_364_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_364_update_start_
      -- 
    req_1249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(306), ack => W_fetch_val3_332_delayed_13_0_362_inst_req_1); -- 
    access_T_cp_element_group_306: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_306"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(308);
      gj_access_T_cp_element_group_306 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(306), clk => clk, reset => reset); --
    end block;
    -- CP-element group 307:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: successors 
    -- CP-element group 307: marked-successors 
    -- CP-element group 307: 	147 
    -- CP-element group 307: 	305 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_364_Sample/ack
      -- CP-element group 307: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_364_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_364_Sample/$exit
      -- 
    ack_1245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val3_332_delayed_13_0_362_inst_ack_0, ack => access_T_CP_0_elements(307)); -- 
    -- CP-element group 308:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	306 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	313 
    -- CP-element group 308: marked-successors 
    -- CP-element group 308: 	146 
    -- CP-element group 308: 	306 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_364_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_364_Update/ack
      -- CP-element group 308: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/assign_stmt_364_Update/$exit
      -- 
    ack_1250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val3_332_delayed_13_0_362_inst_ack_1, ack => access_T_CP_0_elements(308)); -- 
    -- CP-element group 309:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	75 
    -- CP-element group 309: 	151 
    -- CP-element group 309: 	170 
    -- CP-element group 309: marked-predecessors 
    -- CP-element group 309: 	311 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe3_372_sample_start_
      -- CP-element group 309: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe3_372_Sample/$entry
      -- CP-element group 309: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe3_372_Sample/req
      -- 
    req_1258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(309), ack => WPIPE_input_pipe3_372_inst_req_0); -- 
    access_T_cp_element_group_309: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_309"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(75) & access_T_CP_0_elements(151) & access_T_CP_0_elements(170) & access_T_CP_0_elements(311);
      gj_access_T_cp_element_group_309 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(309), clk => clk, reset => reset); --
    end block;
    -- CP-element group 310:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310: marked-successors 
    -- CP-element group 310: 	71 
    -- CP-element group 310: 	147 
    -- CP-element group 310: 	166 
    -- CP-element group 310:  members (6) 
      -- CP-element group 310: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe3_372_sample_completed_
      -- CP-element group 310: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe3_372_update_start_
      -- CP-element group 310: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe3_372_Sample/$exit
      -- CP-element group 310: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe3_372_Sample/ack
      -- CP-element group 310: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe3_372_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe3_372_Update/req
      -- 
    ack_1259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe3_372_inst_ack_0, ack => access_T_CP_0_elements(310)); -- 
    req_1263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(310), ack => WPIPE_input_pipe3_372_inst_req_1); -- 
    -- CP-element group 311:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	313 
    -- CP-element group 311: marked-successors 
    -- CP-element group 311: 	309 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe3_372_update_completed_
      -- CP-element group 311: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe3_372_Update/$exit
      -- CP-element group 311: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/WPIPE_input_pipe3_372_Update/ack
      -- 
    ack_1264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe3_372_inst_ack_1, ack => access_T_CP_0_elements(311)); -- 
    -- CP-element group 312:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	24 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	25 
    -- CP-element group 312:  members (1) 
      -- CP-element group 312: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group access_T_CP_0_elements(312) is a control-delay.
    cp_element_312_delay: control_delay_element  generic map(name => " 312_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(24), ack => access_T_CP_0_elements(312), clk => clk, reset =>reset);
    -- CP-element group 313:  join  transition  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	27 
    -- CP-element group 313: 	229 
    -- CP-element group 313: 	240 
    -- CP-element group 313: 	244 
    -- CP-element group 313: 	248 
    -- CP-element group 313: 	251 
    -- CP-element group 313: 	259 
    -- CP-element group 313: 	270 
    -- CP-element group 313: 	274 
    -- CP-element group 313: 	278 
    -- CP-element group 313: 	281 
    -- CP-element group 313: 	289 
    -- CP-element group 313: 	300 
    -- CP-element group 313: 	304 
    -- CP-element group 313: 	308 
    -- CP-element group 313: 	311 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	21 
    -- CP-element group 313:  members (1) 
      -- CP-element group 313: 	 branch_block_stmt_26/do_while_stmt_79/do_while_stmt_79_loop_body/$exit
      -- 
    access_T_cp_element_group_313: block -- 
      constant place_capacities: IntegerArray(0 to 15) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15);
      constant place_markings: IntegerArray(0 to 15)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant place_delays: IntegerArray(0 to 15) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_313"; 
      signal preds: BooleanArray(1 to 16); -- 
    begin -- 
      preds <= access_T_CP_0_elements(27) & access_T_CP_0_elements(229) & access_T_CP_0_elements(240) & access_T_CP_0_elements(244) & access_T_CP_0_elements(248) & access_T_CP_0_elements(251) & access_T_CP_0_elements(259) & access_T_CP_0_elements(270) & access_T_CP_0_elements(274) & access_T_CP_0_elements(278) & access_T_CP_0_elements(281) & access_T_CP_0_elements(289) & access_T_CP_0_elements(300) & access_T_CP_0_elements(304) & access_T_CP_0_elements(308) & access_T_CP_0_elements(311);
      gj_access_T_cp_element_group_313 : generic_join generic map(name => joinName, number_of_predecessors => 16, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(313), clk => clk, reset => reset); --
    end block;
    -- CP-element group 314:  transition  input  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	20 
    -- CP-element group 314: successors 
    -- CP-element group 314:  members (2) 
      -- CP-element group 314: 	 branch_block_stmt_26/do_while_stmt_79/loop_exit/$exit
      -- CP-element group 314: 	 branch_block_stmt_26/do_while_stmt_79/loop_exit/ack
      -- 
    ack_1269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_79_branch_ack_0, ack => access_T_CP_0_elements(314)); -- 
    -- CP-element group 315:  transition  input  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	20 
    -- CP-element group 315: successors 
    -- CP-element group 315:  members (2) 
      -- CP-element group 315: 	 branch_block_stmt_26/do_while_stmt_79/loop_taken/$exit
      -- CP-element group 315: 	 branch_block_stmt_26/do_while_stmt_79/loop_taken/ack
      -- 
    ack_1273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_79_branch_ack_1, ack => access_T_CP_0_elements(315)); -- 
    -- CP-element group 316:  transition  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	18 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	1 
    -- CP-element group 316:  members (1) 
      -- CP-element group 316: 	 branch_block_stmt_26/do_while_stmt_79/$exit
      -- 
    access_T_CP_0_elements(316) <= access_T_CP_0_elements(18);
    access_T_do_while_stmt_79_terminator_1274: loop_terminator -- 
      generic map (name => " access_T_do_while_stmt_79_terminator_1274", max_iterations_in_flight =>15) 
      port map(loop_body_exit => access_T_CP_0_elements(21),loop_continue => access_T_CP_0_elements(315),loop_terminate => access_T_CP_0_elements(314),loop_back => access_T_CP_0_elements(19),loop_exit => access_T_CP_0_elements(18),clk => clk, reset => reset); -- 
    phi_stmt_81_phi_seq_320_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(36);
      access_T_CP_0_elements(41)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(43);
      access_T_CP_0_elements(42)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(44);
      access_T_CP_0_elements(37) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(38);
      access_T_CP_0_elements(45)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(45);
      access_T_CP_0_elements(46)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(47);
      access_T_CP_0_elements(39) <= phi_mux_reqs(1);
      phi_stmt_81_phi_seq_320 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_81_phi_seq_320") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(32), 
          phi_sample_ack => access_T_CP_0_elements(33), 
          phi_update_req => access_T_CP_0_elements(34), 
          phi_update_ack => access_T_CP_0_elements(35), 
          phi_mux_ack => access_T_CP_0_elements(40), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_86_phi_seq_374_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(55);
      access_T_CP_0_elements(60)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(62);
      access_T_CP_0_elements(61)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(63);
      access_T_CP_0_elements(56) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(57);
      access_T_CP_0_elements(64)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(68);
      access_T_CP_0_elements(65)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(69);
      access_T_CP_0_elements(58) <= phi_mux_reqs(1);
      phi_stmt_86_phi_seq_374 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_86_phi_seq_374") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(51), 
          phi_sample_ack => access_T_CP_0_elements(52), 
          phi_update_req => access_T_CP_0_elements(53), 
          phi_update_ack => access_T_CP_0_elements(54), 
          phi_mux_ack => access_T_CP_0_elements(59), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_91_phi_seq_428_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(76);
      access_T_CP_0_elements(81)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(83);
      access_T_CP_0_elements(82)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(84);
      access_T_CP_0_elements(77) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(78);
      access_T_CP_0_elements(85)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(89);
      access_T_CP_0_elements(86)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(90);
      access_T_CP_0_elements(79) <= phi_mux_reqs(1);
      phi_stmt_91_phi_seq_428 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_91_phi_seq_428") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(72), 
          phi_sample_ack => access_T_CP_0_elements(73), 
          phi_update_req => access_T_CP_0_elements(74), 
          phi_update_ack => access_T_CP_0_elements(75), 
          phi_mux_ack => access_T_CP_0_elements(80), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_96_phi_seq_472_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(95);
      access_T_CP_0_elements(100)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(102);
      access_T_CP_0_elements(101)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(103);
      access_T_CP_0_elements(96) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(97);
      access_T_CP_0_elements(104)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(104);
      access_T_CP_0_elements(105)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(106);
      access_T_CP_0_elements(98) <= phi_mux_reqs(1);
      phi_stmt_96_phi_seq_472 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_96_phi_seq_472") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(26), 
          phi_sample_ack => access_T_CP_0_elements(93), 
          phi_update_req => access_T_CP_0_elements(28), 
          phi_update_ack => access_T_CP_0_elements(94), 
          phi_mux_ack => access_T_CP_0_elements(99), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_101_phi_seq_526_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(114);
      access_T_CP_0_elements(119)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(121);
      access_T_CP_0_elements(120)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(122);
      access_T_CP_0_elements(115) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(116);
      access_T_CP_0_elements(123)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(125);
      access_T_CP_0_elements(124)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(126);
      access_T_CP_0_elements(117) <= phi_mux_reqs(1);
      phi_stmt_101_phi_seq_526 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_101_phi_seq_526") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(110), 
          phi_sample_ack => access_T_CP_0_elements(111), 
          phi_update_req => access_T_CP_0_elements(112), 
          phi_update_ack => access_T_CP_0_elements(113), 
          phi_mux_ack => access_T_CP_0_elements(118), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_105_phi_seq_580_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(133);
      access_T_CP_0_elements(138)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(140);
      access_T_CP_0_elements(139)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(141);
      access_T_CP_0_elements(134) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(135);
      access_T_CP_0_elements(142)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(144);
      access_T_CP_0_elements(143)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(145);
      access_T_CP_0_elements(136) <= phi_mux_reqs(1);
      phi_stmt_105_phi_seq_580 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_105_phi_seq_580") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(129), 
          phi_sample_ack => access_T_CP_0_elements(130), 
          phi_update_req => access_T_CP_0_elements(131), 
          phi_update_ack => access_T_CP_0_elements(132), 
          phi_mux_ack => access_T_CP_0_elements(137), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_109_phi_seq_634_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(152);
      access_T_CP_0_elements(157)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(159);
      access_T_CP_0_elements(158)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(160);
      access_T_CP_0_elements(153) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(154);
      access_T_CP_0_elements(161)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(163);
      access_T_CP_0_elements(162)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(164);
      access_T_CP_0_elements(155) <= phi_mux_reqs(1);
      phi_stmt_109_phi_seq_634 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_109_phi_seq_634") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(148), 
          phi_sample_ack => access_T_CP_0_elements(149), 
          phi_update_req => access_T_CP_0_elements(150), 
          phi_update_ack => access_T_CP_0_elements(151), 
          phi_mux_ack => access_T_CP_0_elements(156), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_113_phi_seq_678_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(171);
      access_T_CP_0_elements(176)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(178);
      access_T_CP_0_elements(177)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(179);
      access_T_CP_0_elements(172) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(173);
      access_T_CP_0_elements(180)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(180);
      access_T_CP_0_elements(181)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(182);
      access_T_CP_0_elements(174) <= phi_mux_reqs(1);
      phi_stmt_113_phi_seq_678 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_113_phi_seq_678") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(167), 
          phi_sample_ack => access_T_CP_0_elements(168), 
          phi_update_req => access_T_CP_0_elements(169), 
          phi_update_ack => access_T_CP_0_elements(170), 
          phi_mux_ack => access_T_CP_0_elements(175), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_118_phi_seq_722_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(192);
      access_T_CP_0_elements(195)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(195);
      access_T_CP_0_elements(196)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(197);
      access_T_CP_0_elements(193) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(190);
      access_T_CP_0_elements(199)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(201);
      access_T_CP_0_elements(200)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(202);
      access_T_CP_0_elements(191) <= phi_mux_reqs(1);
      phi_stmt_118_phi_seq_722 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_118_phi_seq_722") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(186), 
          phi_sample_ack => access_T_CP_0_elements(187), 
          phi_update_req => access_T_CP_0_elements(188), 
          phi_update_ack => access_T_CP_0_elements(189), 
          phi_mux_ack => access_T_CP_0_elements(194), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_123_phi_seq_766_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(211);
      access_T_CP_0_elements(214)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(214);
      access_T_CP_0_elements(215)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(216);
      access_T_CP_0_elements(212) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(209);
      access_T_CP_0_elements(218)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(220);
      access_T_CP_0_elements(219)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(221);
      access_T_CP_0_elements(210) <= phi_mux_reqs(1);
      phi_stmt_123_phi_seq_766 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_123_phi_seq_766") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(205), 
          phi_sample_ack => access_T_CP_0_elements(206), 
          phi_update_req => access_T_CP_0_elements(207), 
          phi_update_ack => access_T_CP_0_elements(208), 
          phi_mux_ack => access_T_CP_0_elements(213), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_272_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= access_T_CP_0_elements(22);
        preds(1)  <= access_T_CP_0_elements(23);
        entry_tmerge_272 : transition_merge -- 
          generic map(name => " entry_tmerge_272")
          port map (preds => preds, symbol_out => access_T_CP_0_elements(24));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_166_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_240_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_314_wire : std_logic_vector(15 downto 0);
    signal ADD_u32_u32_139_wire : std_logic_vector(31 downto 0);
    signal AND_u64_u64_151_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_225_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_299_wire : std_logic_vector(63 downto 0);
    signal LSHR_u32_u32_56_wire : std_logic_vector(31 downto 0);
    signal LSHR_u32_u32_70_wire : std_logic_vector(31 downto 0);
    signal LSHR_u64_u64_159_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_181_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_184_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_194_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_194_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_194_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_233_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_255_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_258_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_268_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_268_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_268_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_307_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_329_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_332_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_347_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_347_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_347_wire : std_logic_vector(63 downto 0);
    signal MUL_u16_u16_31_wire : std_logic_vector(15 downto 0);
    signal NEQ_u64_u1_185_wire : std_logic_vector(0 downto 0);
    signal NEQ_u64_u1_259_wire : std_logic_vector(0 downto 0);
    signal NEQ_u64_u1_333_wire : std_logic_vector(0 downto 0);
    signal SUB_u64_u64_152_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_226_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_300_wire : std_logic_vector(63 downto 0);
    signal address1_81 : std_logic_vector(63 downto 0);
    signal address2_86 : std_logic_vector(63 downto 0);
    signal address3_91 : std_logic_vector(63 downto 0);
    signal array_obj_ref_195_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_195_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_195_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_195_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_195_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_195_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_269_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_269_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_269_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_269_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_269_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_269_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_348_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_348_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_348_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_348_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_348_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_348_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_58_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_58_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_58_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_58_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_58_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_58_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_72_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_72_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_72_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_72_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_72_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_72_root_address : std_logic_vector(13 downto 0);
    signal continue_146 : std_logic_vector(0 downto 0);
    signal continue_183_delayed_1_0_177 : std_logic_vector(0 downto 0);
    signal continue_245_delayed_1_0_251 : std_logic_vector(0 downto 0);
    signal continue_307_delayed_1_0_325 : std_logic_vector(0 downto 0);
    signal fetch_add1_46 : std_logic_vector(31 downto 0);
    signal fetch_add2_60 : std_logic_vector(31 downto 0);
    signal fetch_add3_74 : std_logic_vector(31 downto 0);
    signal fetch_addr1_197 : std_logic_vector(31 downto 0);
    signal fetch_addr2_271 : std_logic_vector(31 downto 0);
    signal fetch_addr3_350 : std_logic_vector(31 downto 0);
    signal fetch_val1_101 : std_logic_vector(63 downto 0);
    signal fetch_val1_203_delayed_13_0_211 : std_logic_vector(63 downto 0);
    signal fetch_val2_105 : std_logic_vector(63 downto 0);
    signal fetch_val2_265_delayed_13_0_285 : std_logic_vector(63 downto 0);
    signal fetch_val3_109 : std_logic_vector(63 downto 0);
    signal fetch_val3_332_delayed_13_0_364 : std_logic_vector(63 downto 0);
    signal fn1_188 : std_logic_vector(0 downto 0);
    signal fn1_195_delayed_7_0_200 : std_logic_vector(0 downto 0);
    signal fn1_201_delayed_13_0_208 : std_logic_vector(0 downto 0);
    signal fn2_257_delayed_7_0_274 : std_logic_vector(0 downto 0);
    signal fn2_262 : std_logic_vector(0 downto 0);
    signal fn2_263_delayed_13_0_282 : std_logic_vector(0 downto 0);
    signal fn3_324_delayed_7_0_353 : std_logic_vector(0 downto 0);
    signal fn3_330_delayed_13_0_361 : std_logic_vector(0 downto 0);
    signal fn3_336 : std_logic_vector(0 downto 0);
    signal fv1_205 : std_logic_vector(63 downto 0);
    signal fv2_279 : std_logic_vector(63 downto 0);
    signal fv3_358 : std_logic_vector(63 downto 0);
    signal konst_136_wire_constant : std_logic_vector(31 downto 0);
    signal konst_138_wire_constant : std_logic_vector(31 downto 0);
    signal konst_148_wire_constant : std_logic_vector(63 downto 0);
    signal konst_150_wire_constant : std_logic_vector(63 downto 0);
    signal konst_153_wire_constant : std_logic_vector(63 downto 0);
    signal konst_165_wire_constant : std_logic_vector(15 downto 0);
    signal konst_172_wire_constant : std_logic_vector(63 downto 0);
    signal konst_180_wire_constant : std_logic_vector(63 downto 0);
    signal konst_183_wire_constant : std_logic_vector(63 downto 0);
    signal konst_193_wire_constant : std_logic_vector(63 downto 0);
    signal konst_222_wire_constant : std_logic_vector(63 downto 0);
    signal konst_224_wire_constant : std_logic_vector(63 downto 0);
    signal konst_227_wire_constant : std_logic_vector(63 downto 0);
    signal konst_239_wire_constant : std_logic_vector(15 downto 0);
    signal konst_246_wire_constant : std_logic_vector(63 downto 0);
    signal konst_254_wire_constant : std_logic_vector(63 downto 0);
    signal konst_257_wire_constant : std_logic_vector(63 downto 0);
    signal konst_267_wire_constant : std_logic_vector(63 downto 0);
    signal konst_296_wire_constant : std_logic_vector(63 downto 0);
    signal konst_298_wire_constant : std_logic_vector(63 downto 0);
    signal konst_301_wire_constant : std_logic_vector(63 downto 0);
    signal konst_313_wire_constant : std_logic_vector(15 downto 0);
    signal konst_320_wire_constant : std_logic_vector(63 downto 0);
    signal konst_328_wire_constant : std_logic_vector(63 downto 0);
    signal konst_331_wire_constant : std_logic_vector(63 downto 0);
    signal konst_346_wire_constant : std_logic_vector(63 downto 0);
    signal konst_36_wire_constant : std_logic_vector(31 downto 0);
    signal konst_55_wire_constant : std_logic_vector(31 downto 0);
    signal konst_69_wire_constant : std_logic_vector(31 downto 0);
    signal m2_factor_38 : std_logic_vector(31 downto 0);
    signal m_factor_33 : std_logic_vector(31 downto 0);
    signal my_fetch1_50 : std_logic_vector(63 downto 0);
    signal my_fetch1_50_104_buffered : std_logic_vector(63 downto 0);
    signal my_fetch2_64 : std_logic_vector(63 downto 0);
    signal my_fetch2_64_108_buffered : std_logic_vector(63 downto 0);
    signal my_fetch3_78 : std_logic_vector(63 downto 0);
    signal my_fetch3_78_112_buffered : std_logic_vector(63 downto 0);
    signal my_num1_155 : std_logic_vector(63 downto 0);
    signal my_num2_229 : std_logic_vector(63 downto 0);
    signal my_num3_303 : std_logic_vector(63 downto 0);
    signal mycounter_96 : std_logic_vector(31 downto 0);
    signal n_address1_174 : std_logic_vector(63 downto 0);
    signal n_address1_174_83_buffered : std_logic_vector(63 downto 0);
    signal n_address2_248 : std_logic_vector(63 downto 0);
    signal n_address2_248_88_buffered : std_logic_vector(63 downto 0);
    signal n_address3_322 : std_logic_vector(63 downto 0);
    signal n_address3_322_93_buffered : std_logic_vector(63 downto 0);
    signal n_fetch_val1_217 : std_logic_vector(63 downto 0);
    signal n_fetch_val1_217_103_buffered : std_logic_vector(63 downto 0);
    signal n_fetch_val2_291 : std_logic_vector(63 downto 0);
    signal n_fetch_val2_291_107_buffered : std_logic_vector(63 downto 0);
    signal n_fetch_val3_370 : std_logic_vector(63 downto 0);
    signal n_fetch_val3_370_111_buffered : std_logic_vector(63 downto 0);
    signal n_mycounter_141 : std_logic_vector(31 downto 0);
    signal n_mycounter_141_98_buffered : std_logic_vector(31 downto 0);
    signal n_row1_169 : std_logic_vector(15 downto 0);
    signal n_row1_169_115_buffered : std_logic_vector(15 downto 0);
    signal n_row2_243 : std_logic_vector(15 downto 0);
    signal n_row2_243_122_buffered : std_logic_vector(15 downto 0);
    signal n_row3_317 : std_logic_vector(15 downto 0);
    signal n_row3_317_127_buffered : std_logic_vector(15 downto 0);
    signal next_row_133 : std_logic_vector(0 downto 0);
    signal ptr_deref_204_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_204_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_204_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_204_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_204_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_278_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_278_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_278_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_278_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_278_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_357_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_357_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_357_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_357_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_357_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_49_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_49_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_49_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_49_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_49_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_63_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_63_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_63_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_63_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_63_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_77_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_77_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_77_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_77_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_77_word_offset_0 : std_logic_vector(13 downto 0);
    signal row1_113 : std_logic_vector(15 downto 0);
    signal row2_118 : std_logic_vector(15 downto 0);
    signal row3_123 : std_logic_vector(15 downto 0);
    signal send_now3_341 : std_logic_vector(0 downto 0);
    signal type_cast_100_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_117_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_121_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_126_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_57_resized : std_logic_vector(13 downto 0);
    signal type_cast_57_scaled : std_logic_vector(13 downto 0);
    signal type_cast_57_wire : std_logic_vector(63 downto 0);
    signal type_cast_71_resized : std_logic_vector(13 downto 0);
    signal type_cast_71_scaled : std_logic_vector(13 downto 0);
    signal type_cast_71_wire : std_logic_vector(63 downto 0);
    signal type_cast_85_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_90_wire : std_logic_vector(63 downto 0);
    signal type_cast_95_wire : std_logic_vector(63 downto 0);
    signal var_val1_161 : std_logic_vector(15 downto 0);
    signal var_val2_235 : std_logic_vector(15 downto 0);
    signal var_val3_309 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_195_constant_part_of_offset <= "00000000000000";
    array_obj_ref_195_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_195_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_195_resized_base_address <= "00000000000000";
    array_obj_ref_269_constant_part_of_offset <= "00000000000000";
    array_obj_ref_269_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_269_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_269_resized_base_address <= "00000000000000";
    array_obj_ref_348_constant_part_of_offset <= "00000000000000";
    array_obj_ref_348_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_348_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_348_resized_base_address <= "00000000000000";
    array_obj_ref_58_constant_part_of_offset <= "00000000000000";
    array_obj_ref_58_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_58_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_58_resized_base_address <= "00000000000000";
    array_obj_ref_72_constant_part_of_offset <= "00000000000000";
    array_obj_ref_72_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_72_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_72_resized_base_address <= "00000000000000";
    fetch_add1_46 <= "00000000000000000000000000000000";
    konst_136_wire_constant <= "00000000000000000000000000000001";
    konst_138_wire_constant <= "00000000000000000000000000000001";
    konst_148_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_150_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_153_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_165_wire_constant <= "0000000000000001";
    konst_172_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_180_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_183_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_193_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_222_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_224_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_227_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_239_wire_constant <= "0000000000000001";
    konst_246_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_254_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_257_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_267_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_296_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_298_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_301_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_313_wire_constant <= "0000000000000001";
    konst_320_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_328_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_331_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_346_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_36_wire_constant <= "00000000000000000000000000000001";
    konst_55_wire_constant <= "00000000000000000000000000000010";
    konst_69_wire_constant <= "00000000000000000000000000000001";
    ptr_deref_204_word_offset_0 <= "00000000000000";
    ptr_deref_278_word_offset_0 <= "00000000000000";
    ptr_deref_357_word_offset_0 <= "00000000000000";
    ptr_deref_49_word_offset_0 <= "00000000000000";
    ptr_deref_63_word_offset_0 <= "00000000000000";
    ptr_deref_77_word_offset_0 <= "00000000000000";
    type_cast_100_wire_constant <= "00000000000000000000000000000001";
    type_cast_117_wire_constant <= "0000000000000000";
    type_cast_121_wire_constant <= "0000000000000001";
    type_cast_126_wire_constant <= "0000000000000010";
    type_cast_85_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_101: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_fetch_val1_217_103_buffered & my_fetch1_50_104_buffered;
      req <= phi_stmt_101_req_0 & phi_stmt_101_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_101",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_101_ack_0,
          idata => idata,
          odata => fetch_val1_101,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_101
    phi_stmt_105: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_fetch_val2_291_107_buffered & my_fetch2_64_108_buffered;
      req <= phi_stmt_105_req_0 & phi_stmt_105_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_105",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_105_ack_0,
          idata => idata,
          odata => fetch_val2_105,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_105
    phi_stmt_109: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_fetch_val3_370_111_buffered & my_fetch3_78_112_buffered;
      req <= phi_stmt_109_req_0 & phi_stmt_109_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_109",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_109_ack_0,
          idata => idata,
          odata => fetch_val3_109,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_109
    phi_stmt_113: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_row1_169_115_buffered & type_cast_117_wire_constant;
      req <= phi_stmt_113_req_0 & phi_stmt_113_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_113",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_113_ack_0,
          idata => idata,
          odata => row1_113,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_113
    phi_stmt_118: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_121_wire_constant & n_row2_243_122_buffered;
      req <= phi_stmt_118_req_0 & phi_stmt_118_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_118",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_118_ack_0,
          idata => idata,
          odata => row2_118,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_118
    phi_stmt_123: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_126_wire_constant & n_row3_317_127_buffered;
      req <= phi_stmt_123_req_0 & phi_stmt_123_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_123",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_123_ack_0,
          idata => idata,
          odata => row3_123,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_123
    phi_stmt_81: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_address1_174_83_buffered & type_cast_85_wire_constant;
      req <= phi_stmt_81_req_0 & phi_stmt_81_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_81",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_81_ack_0,
          idata => idata,
          odata => address1_81,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_81
    phi_stmt_86: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_address2_248_88_buffered & type_cast_90_wire;
      req <= phi_stmt_86_req_0 & phi_stmt_86_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_86",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_86_ack_0,
          idata => idata,
          odata => address2_86,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_86
    phi_stmt_91: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_address3_322_93_buffered & type_cast_95_wire;
      req <= phi_stmt_91_req_0 & phi_stmt_91_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_91",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_91_ack_0,
          idata => idata,
          odata => address3_91,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_91
    phi_stmt_96: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_mycounter_141_98_buffered & type_cast_100_wire_constant;
      req <= phi_stmt_96_req_0 & phi_stmt_96_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_96",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_96_ack_0,
          idata => idata,
          odata => mycounter_96,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_96
    -- flow-through select operator MUX_140_inst
    n_mycounter_141 <= konst_136_wire_constant when (next_row_133(0) /=  '0') else ADD_u32_u32_139_wire;
    -- flow-through select operator MUX_168_inst
    n_row1_169 <= ADD_u16_u16_166_wire when (next_row_133(0) /=  '0') else row1_113;
    -- flow-through select operator MUX_216_inst
    n_fetch_val1_217 <= fv1_205 when (fn1_201_delayed_13_0_208(0) /=  '0') else fetch_val1_203_delayed_13_0_211;
    -- flow-through select operator MUX_242_inst
    n_row2_243 <= ADD_u16_u16_240_wire when (next_row_133(0) /=  '0') else row2_118;
    -- flow-through select operator MUX_290_inst
    n_fetch_val2_291 <= fv2_279 when (fn2_263_delayed_13_0_282(0) /=  '0') else fetch_val2_265_delayed_13_0_285;
    -- flow-through select operator MUX_316_inst
    n_row3_317 <= ADD_u16_u16_314_wire when (next_row_133(0) /=  '0') else row3_123;
    -- flow-through select operator MUX_369_inst
    n_fetch_val3_370 <= fv3_358 when (fn3_330_delayed_13_0_361(0) /=  '0') else fetch_val3_332_delayed_13_0_364;
    W_continue_183_delayed_1_0_175_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_continue_183_delayed_1_0_175_inst_req_0;
      W_continue_183_delayed_1_0_175_inst_ack_0<= wack(0);
      rreq(0) <= W_continue_183_delayed_1_0_175_inst_req_1;
      W_continue_183_delayed_1_0_175_inst_ack_1<= rack(0);
      W_continue_183_delayed_1_0_175_inst : InterlockBuffer generic map ( -- 
        name => "W_continue_183_delayed_1_0_175_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => continue_146,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => continue_183_delayed_1_0_177,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_continue_245_delayed_1_0_249_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_continue_245_delayed_1_0_249_inst_req_0;
      W_continue_245_delayed_1_0_249_inst_ack_0<= wack(0);
      rreq(0) <= W_continue_245_delayed_1_0_249_inst_req_1;
      W_continue_245_delayed_1_0_249_inst_ack_1<= rack(0);
      W_continue_245_delayed_1_0_249_inst : InterlockBuffer generic map ( -- 
        name => "W_continue_245_delayed_1_0_249_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => continue_146,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => continue_245_delayed_1_0_251,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_continue_307_delayed_1_0_323_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_continue_307_delayed_1_0_323_inst_req_0;
      W_continue_307_delayed_1_0_323_inst_ack_0<= wack(0);
      rreq(0) <= W_continue_307_delayed_1_0_323_inst_req_1;
      W_continue_307_delayed_1_0_323_inst_ack_1<= rack(0);
      W_continue_307_delayed_1_0_323_inst : InterlockBuffer generic map ( -- 
        name => "W_continue_307_delayed_1_0_323_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => continue_146,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => continue_307_delayed_1_0_325,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fetch_val1_203_delayed_13_0_209_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val1_203_delayed_13_0_209_inst_req_0;
      W_fetch_val1_203_delayed_13_0_209_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val1_203_delayed_13_0_209_inst_req_1;
      W_fetch_val1_203_delayed_13_0_209_inst_ack_1<= rack(0);
      W_fetch_val1_203_delayed_13_0_209_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val1_203_delayed_13_0_209_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val1_101,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val1_203_delayed_13_0_211,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fetch_val2_265_delayed_13_0_283_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val2_265_delayed_13_0_283_inst_req_0;
      W_fetch_val2_265_delayed_13_0_283_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val2_265_delayed_13_0_283_inst_req_1;
      W_fetch_val2_265_delayed_13_0_283_inst_ack_1<= rack(0);
      W_fetch_val2_265_delayed_13_0_283_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val2_265_delayed_13_0_283_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val2_105,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val2_265_delayed_13_0_285,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fetch_val3_332_delayed_13_0_362_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val3_332_delayed_13_0_362_inst_req_0;
      W_fetch_val3_332_delayed_13_0_362_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val3_332_delayed_13_0_362_inst_req_1;
      W_fetch_val3_332_delayed_13_0_362_inst_ack_1<= rack(0);
      W_fetch_val3_332_delayed_13_0_362_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val3_332_delayed_13_0_362_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val3_109,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val3_332_delayed_13_0_364,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn1_195_delayed_7_0_198_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn1_195_delayed_7_0_198_inst_req_0;
      W_fn1_195_delayed_7_0_198_inst_ack_0<= wack(0);
      rreq(0) <= W_fn1_195_delayed_7_0_198_inst_req_1;
      W_fn1_195_delayed_7_0_198_inst_ack_1<= rack(0);
      W_fn1_195_delayed_7_0_198_inst : InterlockBuffer generic map ( -- 
        name => "W_fn1_195_delayed_7_0_198_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn1_188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn1_195_delayed_7_0_200,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn1_201_delayed_13_0_206_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn1_201_delayed_13_0_206_inst_req_0;
      W_fn1_201_delayed_13_0_206_inst_ack_0<= wack(0);
      rreq(0) <= W_fn1_201_delayed_13_0_206_inst_req_1;
      W_fn1_201_delayed_13_0_206_inst_ack_1<= rack(0);
      W_fn1_201_delayed_13_0_206_inst : InterlockBuffer generic map ( -- 
        name => "W_fn1_201_delayed_13_0_206_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn1_188,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn1_201_delayed_13_0_208,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn2_257_delayed_7_0_272_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn2_257_delayed_7_0_272_inst_req_0;
      W_fn2_257_delayed_7_0_272_inst_ack_0<= wack(0);
      rreq(0) <= W_fn2_257_delayed_7_0_272_inst_req_1;
      W_fn2_257_delayed_7_0_272_inst_ack_1<= rack(0);
      W_fn2_257_delayed_7_0_272_inst : InterlockBuffer generic map ( -- 
        name => "W_fn2_257_delayed_7_0_272_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn2_262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn2_257_delayed_7_0_274,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn2_263_delayed_13_0_280_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn2_263_delayed_13_0_280_inst_req_0;
      W_fn2_263_delayed_13_0_280_inst_ack_0<= wack(0);
      rreq(0) <= W_fn2_263_delayed_13_0_280_inst_req_1;
      W_fn2_263_delayed_13_0_280_inst_ack_1<= rack(0);
      W_fn2_263_delayed_13_0_280_inst : InterlockBuffer generic map ( -- 
        name => "W_fn2_263_delayed_13_0_280_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn2_262,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn2_263_delayed_13_0_282,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn3_324_delayed_7_0_351_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn3_324_delayed_7_0_351_inst_req_0;
      W_fn3_324_delayed_7_0_351_inst_ack_0<= wack(0);
      rreq(0) <= W_fn3_324_delayed_7_0_351_inst_req_1;
      W_fn3_324_delayed_7_0_351_inst_ack_1<= rack(0);
      W_fn3_324_delayed_7_0_351_inst : InterlockBuffer generic map ( -- 
        name => "W_fn3_324_delayed_7_0_351_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn3_336,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn3_324_delayed_7_0_353,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn3_330_delayed_13_0_359_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn3_330_delayed_13_0_359_inst_req_0;
      W_fn3_330_delayed_13_0_359_inst_ack_0<= wack(0);
      rreq(0) <= W_fn3_330_delayed_13_0_359_inst_req_1;
      W_fn3_330_delayed_13_0_359_inst_ack_1<= rack(0);
      W_fn3_330_delayed_13_0_359_inst : InterlockBuffer generic map ( -- 
        name => "W_fn3_330_delayed_13_0_359_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn3_336,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn3_330_delayed_13_0_361,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_196_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_196_final_reg_req_0;
      addr_of_196_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_196_final_reg_req_1;
      addr_of_196_final_reg_ack_1<= rack(0);
      addr_of_196_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_196_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_195_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr1_197,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_270_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_270_final_reg_req_0;
      addr_of_270_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_270_final_reg_req_1;
      addr_of_270_final_reg_ack_1<= rack(0);
      addr_of_270_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_270_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_269_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr2_271,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_349_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_349_final_reg_req_0;
      addr_of_349_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_349_final_reg_req_1;
      addr_of_349_final_reg_ack_1<= rack(0);
      addr_of_349_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_349_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_348_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr3_350,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_59_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_59_final_reg_req_0;
      addr_of_59_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_59_final_reg_req_1;
      addr_of_59_final_reg_ack_1<= rack(0);
      addr_of_59_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_59_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_58_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_add2_60,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_73_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_73_final_reg_req_0;
      addr_of_73_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_73_final_reg_req_1;
      addr_of_73_final_reg_ack_1<= rack(0);
      addr_of_73_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_73_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_72_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_add3_74,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch1_50_104_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch1_50_104_buf_req_0;
      my_fetch1_50_104_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch1_50_104_buf_req_1;
      my_fetch1_50_104_buf_ack_1<= rack(0);
      my_fetch1_50_104_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch1_50_104_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch1_50,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch1_50_104_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch2_64_108_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch2_64_108_buf_req_0;
      my_fetch2_64_108_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch2_64_108_buf_req_1;
      my_fetch2_64_108_buf_ack_1<= rack(0);
      my_fetch2_64_108_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch2_64_108_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch2_64,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch2_64_108_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch3_78_112_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch3_78_112_buf_req_0;
      my_fetch3_78_112_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch3_78_112_buf_req_1;
      my_fetch3_78_112_buf_ack_1<= rack(0);
      my_fetch3_78_112_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch3_78_112_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch3_78,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch3_78_112_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address1_174_83_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address1_174_83_buf_req_0;
      n_address1_174_83_buf_ack_0<= wack(0);
      rreq(0) <= n_address1_174_83_buf_req_1;
      n_address1_174_83_buf_ack_1<= rack(0);
      n_address1_174_83_buf : InterlockBuffer generic map ( -- 
        name => "n_address1_174_83_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address1_174,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address1_174_83_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address2_248_88_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address2_248_88_buf_req_0;
      n_address2_248_88_buf_ack_0<= wack(0);
      rreq(0) <= n_address2_248_88_buf_req_1;
      n_address2_248_88_buf_ack_1<= rack(0);
      n_address2_248_88_buf : InterlockBuffer generic map ( -- 
        name => "n_address2_248_88_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address2_248,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address2_248_88_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address3_322_93_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address3_322_93_buf_req_0;
      n_address3_322_93_buf_ack_0<= wack(0);
      rreq(0) <= n_address3_322_93_buf_req_1;
      n_address3_322_93_buf_ack_1<= rack(0);
      n_address3_322_93_buf : InterlockBuffer generic map ( -- 
        name => "n_address3_322_93_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address3_322,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address3_322_93_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_fetch_val1_217_103_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_fetch_val1_217_103_buf_req_0;
      n_fetch_val1_217_103_buf_ack_0<= wack(0);
      rreq(0) <= n_fetch_val1_217_103_buf_req_1;
      n_fetch_val1_217_103_buf_ack_1<= rack(0);
      n_fetch_val1_217_103_buf : InterlockBuffer generic map ( -- 
        name => "n_fetch_val1_217_103_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_fetch_val1_217,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_fetch_val1_217_103_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_fetch_val2_291_107_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_fetch_val2_291_107_buf_req_0;
      n_fetch_val2_291_107_buf_ack_0<= wack(0);
      rreq(0) <= n_fetch_val2_291_107_buf_req_1;
      n_fetch_val2_291_107_buf_ack_1<= rack(0);
      n_fetch_val2_291_107_buf : InterlockBuffer generic map ( -- 
        name => "n_fetch_val2_291_107_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_fetch_val2_291,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_fetch_val2_291_107_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_fetch_val3_370_111_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_fetch_val3_370_111_buf_req_0;
      n_fetch_val3_370_111_buf_ack_0<= wack(0);
      rreq(0) <= n_fetch_val3_370_111_buf_req_1;
      n_fetch_val3_370_111_buf_ack_1<= rack(0);
      n_fetch_val3_370_111_buf : InterlockBuffer generic map ( -- 
        name => "n_fetch_val3_370_111_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_fetch_val3_370,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_fetch_val3_370_111_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_mycounter_141_98_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_mycounter_141_98_buf_req_0;
      n_mycounter_141_98_buf_ack_0<= wack(0);
      rreq(0) <= n_mycounter_141_98_buf_req_1;
      n_mycounter_141_98_buf_ack_1<= rack(0);
      n_mycounter_141_98_buf : InterlockBuffer generic map ( -- 
        name => "n_mycounter_141_98_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_mycounter_141,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_mycounter_141_98_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row1_169_115_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row1_169_115_buf_req_0;
      n_row1_169_115_buf_ack_0<= wack(0);
      rreq(0) <= n_row1_169_115_buf_req_1;
      n_row1_169_115_buf_ack_1<= rack(0);
      n_row1_169_115_buf : InterlockBuffer generic map ( -- 
        name => "n_row1_169_115_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row1_169,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row1_169_115_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row2_243_122_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row2_243_122_buf_req_0;
      n_row2_243_122_buf_ack_0<= wack(0);
      rreq(0) <= n_row2_243_122_buf_req_1;
      n_row2_243_122_buf_ack_1<= rack(0);
      n_row2_243_122_buf : InterlockBuffer generic map ( -- 
        name => "n_row2_243_122_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row2_243,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row2_243_122_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row3_317_127_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row3_317_127_buf_req_0;
      n_row3_317_127_buf_ack_0<= wack(0);
      rreq(0) <= n_row3_317_127_buf_req_1;
      n_row3_317_127_buf_ack_1<= rack(0);
      n_row3_317_127_buf : InterlockBuffer generic map ( -- 
        name => "n_row3_317_127_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row3_317,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row3_317_127_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_160_inst
    process(LSHR_u64_u64_159_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_159_wire(15 downto 0);
      var_val1_161 <= tmp_var; -- 
    end process;
    -- interlock type_cast_234_inst
    process(LSHR_u64_u64_233_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_233_wire(15 downto 0);
      var_val2_235 <= tmp_var; -- 
    end process;
    -- interlock type_cast_308_inst
    process(LSHR_u64_u64_307_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_307_wire(15 downto 0);
      var_val3_309 <= tmp_var; -- 
    end process;
    -- interlock type_cast_32_inst
    process(MUL_u16_u16_31_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_31_wire(15 downto 0);
      m_factor_33 <= tmp_var; -- 
    end process;
    -- interlock type_cast_57_inst
    process(LSHR_u32_u32_56_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_56_wire(31 downto 0);
      type_cast_57_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_71_inst
    process(LSHR_u32_u32_70_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_70_wire(31 downto 0);
      type_cast_71_wire <= tmp_var; -- 
    end process;
    type_cast_90_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_90_inst_req_0;
      type_cast_90_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_90_inst_req_1;
      type_cast_90_inst_ack_1<= rack(0);
      type_cast_90_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_90_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_33,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_90_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_95_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_95_inst_req_0;
      type_cast_95_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_95_inst_req_1;
      type_cast_95_inst_ack_1<= rack(0);
      type_cast_95_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_95_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m2_factor_38,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_95_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_195_index_1_rename
    process(LSHR_u64_u64_194_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_194_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_194_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_195_index_1_resize
    process(LSHR_u64_u64_194_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_194_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_194_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_195_root_address_inst
    process(array_obj_ref_195_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_195_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_195_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_269_index_1_rename
    process(LSHR_u64_u64_268_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_268_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_268_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_269_index_1_resize
    process(LSHR_u64_u64_268_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_268_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_268_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_269_root_address_inst
    process(array_obj_ref_269_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_269_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_269_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_348_index_1_rename
    process(LSHR_u64_u64_347_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_347_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_347_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_348_index_1_resize
    process(LSHR_u64_u64_347_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_347_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_347_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_348_root_address_inst
    process(array_obj_ref_348_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_348_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_348_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_58_index_1_rename
    process(type_cast_57_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_57_resized;
      ov(13 downto 0) := iv;
      type_cast_57_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_58_index_1_resize
    process(type_cast_57_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_57_wire;
      ov := iv(13 downto 0);
      type_cast_57_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_58_root_address_inst
    process(array_obj_ref_58_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_58_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_58_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_72_index_1_rename
    process(type_cast_71_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_71_resized;
      ov(13 downto 0) := iv;
      type_cast_71_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_72_index_1_resize
    process(type_cast_71_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_71_wire;
      ov := iv(13 downto 0);
      type_cast_71_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_72_root_address_inst
    process(array_obj_ref_72_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_72_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_72_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_204_addr_0
    process(ptr_deref_204_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_204_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_204_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_204_base_resize
    process(fetch_addr1_197) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr1_197;
      ov := iv(13 downto 0);
      ptr_deref_204_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_204_gather_scatter
    process(ptr_deref_204_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_204_data_0;
      ov(63 downto 0) := iv;
      fv1_205 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_204_root_address_inst
    process(ptr_deref_204_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_204_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_204_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_278_addr_0
    process(ptr_deref_278_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_278_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_278_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_278_base_resize
    process(fetch_addr2_271) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr2_271;
      ov := iv(13 downto 0);
      ptr_deref_278_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_278_gather_scatter
    process(ptr_deref_278_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_278_data_0;
      ov(63 downto 0) := iv;
      fv2_279 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_278_root_address_inst
    process(ptr_deref_278_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_278_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_278_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_357_addr_0
    process(ptr_deref_357_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_357_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_357_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_357_base_resize
    process(fetch_addr3_350) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr3_350;
      ov := iv(13 downto 0);
      ptr_deref_357_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_357_gather_scatter
    process(ptr_deref_357_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_357_data_0;
      ov(63 downto 0) := iv;
      fv3_358 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_357_root_address_inst
    process(ptr_deref_357_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_357_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_357_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_49_addr_0
    process(ptr_deref_49_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_49_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_49_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_49_base_resize
    process(fetch_add1_46) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_add1_46;
      ov := iv(13 downto 0);
      ptr_deref_49_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_49_gather_scatter
    process(ptr_deref_49_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_49_data_0;
      ov(63 downto 0) := iv;
      my_fetch1_50 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_49_root_address_inst
    process(ptr_deref_49_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_49_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_49_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_63_addr_0
    process(ptr_deref_63_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_63_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_63_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_63_base_resize
    process(fetch_add2_60) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_add2_60;
      ov := iv(13 downto 0);
      ptr_deref_63_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_63_gather_scatter
    process(ptr_deref_63_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_63_data_0;
      ov(63 downto 0) := iv;
      my_fetch2_64 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_63_root_address_inst
    process(ptr_deref_63_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_63_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_63_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_77_addr_0
    process(ptr_deref_77_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_77_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_77_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_77_base_resize
    process(fetch_add3_74) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_add3_74;
      ov := iv(13 downto 0);
      ptr_deref_77_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_77_gather_scatter
    process(ptr_deref_77_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_77_data_0;
      ov(63 downto 0) := iv;
      my_fetch3_78 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_77_root_address_inst
    process(ptr_deref_77_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_77_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_77_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_79_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_146;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_79_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_79_branch_req_0,
          ack0 => do_while_stmt_79_branch_ack_0,
          ack1 => do_while_stmt_79_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_166_inst
    process(row1_113) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row1_113, konst_165_wire_constant, tmp_var);
      ADD_u16_u16_166_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_240_inst
    process(row2_118) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row2_118, konst_239_wire_constant, tmp_var);
      ADD_u16_u16_240_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_314_inst
    process(row3_123) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row3_123, konst_313_wire_constant, tmp_var);
      ADD_u16_u16_314_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_139_inst
    process(mycounter_96) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycounter_96, konst_138_wire_constant, tmp_var);
      ADD_u32_u32_139_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_173_inst
    process(address1_81) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address1_81, konst_172_wire_constant, tmp_var);
      n_address1_174 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_247_inst
    process(address2_86) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address2_86, konst_246_wire_constant, tmp_var);
      n_address2_248 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_321_inst
    process(address3_91) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address3_91, konst_320_wire_constant, tmp_var);
      n_address3_322 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_187_inst
    process(NEQ_u64_u1_185_wire, continue_183_delayed_1_0_177) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u64_u1_185_wire, continue_183_delayed_1_0_177, tmp_var);
      fn1_188 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_261_inst
    process(NEQ_u64_u1_259_wire, continue_245_delayed_1_0_251) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u64_u1_259_wire, continue_245_delayed_1_0_251, tmp_var);
      fn2_262 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_335_inst
    process(NEQ_u64_u1_333_wire, continue_307_delayed_1_0_325) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u64_u1_333_wire, continue_307_delayed_1_0_325, tmp_var);
      fn3_336 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_151_inst
    process(address1_81) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(address1_81, konst_150_wire_constant, tmp_var);
      AND_u64_u64_151_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_225_inst
    process(address2_86) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(address2_86, konst_224_wire_constant, tmp_var);
      AND_u64_u64_225_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_299_inst
    process(address3_91) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(address3_91, konst_298_wire_constant, tmp_var);
      AND_u64_u64_299_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_132_inst
    process(mycounter_96, m_factor_33) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(mycounter_96, m_factor_33, tmp_var);
      next_row_133 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_56_inst
    process(m_factor_33) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(m_factor_33, konst_55_wire_constant, tmp_var);
      LSHR_u32_u32_56_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_70_inst
    process(m_factor_33) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(m_factor_33, konst_69_wire_constant, tmp_var);
      LSHR_u32_u32_70_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_159_inst
    process(fetch_val1_101, my_num1_155) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val1_101, my_num1_155, tmp_var);
      LSHR_u64_u64_159_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_181_inst
    process(n_address1_174) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address1_174, konst_180_wire_constant, tmp_var);
      LSHR_u64_u64_181_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_184_inst
    process(address1_81) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address1_81, konst_183_wire_constant, tmp_var);
      LSHR_u64_u64_184_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_194_inst
    process(n_address1_174) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address1_174, konst_193_wire_constant, tmp_var);
      LSHR_u64_u64_194_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_233_inst
    process(fetch_val2_105, my_num2_229) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val2_105, my_num2_229, tmp_var);
      LSHR_u64_u64_233_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_255_inst
    process(n_address2_248) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address2_248, konst_254_wire_constant, tmp_var);
      LSHR_u64_u64_255_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_258_inst
    process(address2_86) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address2_86, konst_257_wire_constant, tmp_var);
      LSHR_u64_u64_258_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_268_inst
    process(n_address2_248) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address2_248, konst_267_wire_constant, tmp_var);
      LSHR_u64_u64_268_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_307_inst
    process(fetch_val3_109, my_num3_303) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val3_109, my_num3_303, tmp_var);
      LSHR_u64_u64_307_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_329_inst
    process(n_address3_322) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address3_322, konst_328_wire_constant, tmp_var);
      LSHR_u64_u64_329_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_332_inst
    process(address3_91) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address3_91, konst_331_wire_constant, tmp_var);
      LSHR_u64_u64_332_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_347_inst
    process(n_address3_322) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(n_address3_322, konst_346_wire_constant, tmp_var);
      LSHR_u64_u64_347_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_31_inst
    process(ct_buffer, chl_in_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, chl_in_buffer, tmp_var);
      MUL_u16_u16_31_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u64_u1_185_inst
    process(LSHR_u64_u64_181_wire, LSHR_u64_u64_184_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(LSHR_u64_u64_181_wire, LSHR_u64_u64_184_wire, tmp_var);
      NEQ_u64_u1_185_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u64_u1_259_inst
    process(LSHR_u64_u64_255_wire, LSHR_u64_u64_258_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(LSHR_u64_u64_255_wire, LSHR_u64_u64_258_wire, tmp_var);
      NEQ_u64_u1_259_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u64_u1_333_inst
    process(LSHR_u64_u64_329_wire, LSHR_u64_u64_332_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(LSHR_u64_u64_329_wire, LSHR_u64_u64_332_wire, tmp_var);
      NEQ_u64_u1_333_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_37_inst
    process(m_factor_33) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(m_factor_33, konst_36_wire_constant, tmp_var);
      m2_factor_38 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_154_inst
    process(SUB_u64_u64_152_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_152_wire, konst_153_wire_constant, tmp_var);
      my_num1_155 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_228_inst
    process(SUB_u64_u64_226_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_226_wire, konst_227_wire_constant, tmp_var);
      my_num2_229 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_302_inst
    process(SUB_u64_u64_300_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_300_wire, konst_301_wire_constant, tmp_var);
      my_num3_303 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_152_inst
    process(konst_148_wire_constant, AND_u64_u64_151_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_148_wire_constant, AND_u64_u64_151_wire, tmp_var);
      SUB_u64_u64_152_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_226_inst
    process(konst_222_wire_constant, AND_u64_u64_225_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_222_wire_constant, AND_u64_u64_225_wire, tmp_var);
      SUB_u64_u64_226_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_300_inst
    process(konst_296_wire_constant, AND_u64_u64_299_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_296_wire_constant, AND_u64_u64_299_wire, tmp_var);
      SUB_u64_u64_300_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_145_inst
    process(n_row1_169, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_row1_169, row_in_buffer, tmp_var);
      continue_146 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_340_inst
    process(row1_113, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(row1_113, row_in_buffer, tmp_var);
      send_now3_341 <= tmp_var; --
    end process;
    -- shared split operator group (41) : array_obj_ref_195_index_offset 
    ApIntAdd_group_41: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_194_scaled;
      array_obj_ref_195_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_195_index_offset_req_0;
      array_obj_ref_195_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_195_index_offset_req_1;
      array_obj_ref_195_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_41_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_41_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_41",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : array_obj_ref_269_index_offset 
    ApIntAdd_group_42: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_268_scaled;
      array_obj_ref_269_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_269_index_offset_req_0;
      array_obj_ref_269_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_269_index_offset_req_1;
      array_obj_ref_269_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_42_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_42_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_42",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : array_obj_ref_348_index_offset 
    ApIntAdd_group_43: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_347_scaled;
      array_obj_ref_348_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_348_index_offset_req_0;
      array_obj_ref_348_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_348_index_offset_req_1;
      array_obj_ref_348_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_43_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_43_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_43",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : array_obj_ref_58_index_offset 
    ApIntAdd_group_44: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_57_scaled;
      array_obj_ref_58_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_58_index_offset_req_0;
      array_obj_ref_58_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_58_index_offset_req_1;
      array_obj_ref_58_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_44_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_44_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_44",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : array_obj_ref_72_index_offset 
    ApIntAdd_group_45: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_71_scaled;
      array_obj_ref_72_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_72_index_offset_req_0;
      array_obj_ref_72_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_72_index_offset_req_1;
      array_obj_ref_72_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_45_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_45_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_45",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared load operator group (0) : ptr_deref_63_load_0 ptr_deref_77_load_0 ptr_deref_204_load_0 ptr_deref_49_load_0 ptr_deref_278_load_0 ptr_deref_357_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(83 downto 0);
      signal data_out: std_logic_vector(383 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 5 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 5 downto 0);
      signal guard_vector : std_logic_vector( 5 downto 0);
      constant inBUFs : IntegerArray(5 downto 0) := (5 => 0, 4 => 0, 3 => 2, 2 => 0, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(5 downto 0) := (5 => 1, 4 => 1, 3 => 2, 2 => 1, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(5 downto 0) := (0 => true, 1 => true, 2 => false, 3 => true, 4 => false, 5 => false);
      constant guardBuffering: IntegerArray(5 downto 0)  := (0 => 6, 1 => 6, 2 => 2, 3 => 6, 4 => 2, 5 => 2);
      -- 
    begin -- 
      reqL_unguarded(5) <= ptr_deref_63_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_77_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_204_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_49_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_278_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_357_load_0_req_0;
      ptr_deref_63_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_77_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_204_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_49_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_278_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_357_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(5) <= ptr_deref_63_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_77_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_204_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_49_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_278_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_357_load_0_req_1;
      ptr_deref_63_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_77_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_204_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_49_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_278_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_357_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= fn3_324_delayed_7_0_353(0);
      guard_vector(1)  <= fn2_257_delayed_7_0_274(0);
      guard_vector(2)  <=  '1';
      guard_vector(3)  <= fn1_195_delayed_7_0_200(0);
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 2) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 6, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_63_word_address_0 & ptr_deref_77_word_address_0 & ptr_deref_204_word_address_0 & ptr_deref_49_word_address_0 & ptr_deref_278_word_address_0 & ptr_deref_357_word_address_0;
      ptr_deref_63_data_0 <= data_out(383 downto 320);
      ptr_deref_77_data_0 <= data_out(319 downto 256);
      ptr_deref_204_data_0 <= data_out(255 downto 192);
      ptr_deref_49_data_0 <= data_out(191 downto 128);
      ptr_deref_278_data_0 <= data_out(127 downto 64);
      ptr_deref_357_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 6,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 6,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_input_pipe1_218_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_pipe1_218_inst_req_0;
      WPIPE_input_pipe1_218_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_pipe1_218_inst_req_1;
      WPIPE_input_pipe1_218_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= var_val1_161;
      input_pipe1_write_0_gI: SplitGuardInterface generic map(name => "input_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "input_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe1_pipe_write_req(0),
          oack => input_pipe1_pipe_write_ack(0),
          odata => input_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_input_pipe2_292_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_pipe2_292_inst_req_0;
      WPIPE_input_pipe2_292_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_pipe2_292_inst_req_1;
      WPIPE_input_pipe2_292_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= var_val2_235;
      input_pipe2_write_1_gI: SplitGuardInterface generic map(name => "input_pipe2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe2_write_1: OutputPortRevised -- 
        generic map ( name => "input_pipe2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe2_pipe_write_req(0),
          oack => input_pipe2_pipe_write_ack(0),
          odata => input_pipe2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_input_pipe3_372_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_pipe3_372_inst_req_0;
      WPIPE_input_pipe3_372_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_pipe3_372_inst_req_1;
      WPIPE_input_pipe3_372_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_now3_341(0);
      data_in <= var_val3_309;
      input_pipe3_write_2_gI: SplitGuardInterface generic map(name => "input_pipe3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe3_write_2: OutputPortRevised -- 
        generic map ( name => "input_pipe3", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe3_pipe_write_req(0),
          oack => input_pipe3_pipe_write_ack(0),
          odata => input_pipe3_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- 
  end Block; -- data_path
  -- 
end access_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolution3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    access_T_call_reqs : out  std_logic_vector(0 downto 0);
    access_T_call_acks : in   std_logic_vector(0 downto 0);
    access_T_call_data : out  std_logic_vector(47 downto 0);
    access_T_call_tag  :  out  std_logic_vector(0 downto 0);
    access_T_return_reqs : out  std_logic_vector(0 downto 0);
    access_T_return_acks : in   std_logic_vector(0 downto 0);
    access_T_return_tag :  in   std_logic_vector(0 downto 0);
    loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_call_data : out  std_logic_vector(79 downto 0);
    loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolution3D;
architecture convolution3D_arch of convolution3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolution3D_CP_1767_start: Boolean;
  signal convolution3D_CP_1767_symbol: Boolean;
  -- volatile/operator module components. 
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      row_in : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      input_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      num_chl : in  std_logic_vector(15 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_maxpool_input_pipe_893_inst_ack_0 : boolean;
  signal type_cast_574_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_929_inst_ack_0 : boolean;
  signal array_obj_ref_876_index_offset_req_0 : boolean;
  signal type_cast_884_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_893_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_570_inst_ack_1 : boolean;
  signal type_cast_586_inst_ack_0 : boolean;
  signal type_cast_586_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_929_inst_req_0 : boolean;
  signal ptr_deref_1013_store_0_req_0 : boolean;
  signal type_cast_561_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_929_inst_req_1 : boolean;
  signal type_cast_884_inst_req_0 : boolean;
  signal type_cast_599_inst_ack_1 : boolean;
  signal array_obj_ref_1192_index_offset_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_620_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_620_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1001_inst_req_0 : boolean;
  signal array_obj_ref_876_index_offset_req_1 : boolean;
  signal type_cast_969_inst_req_1 : boolean;
  signal if_stmt_1078_branch_ack_0 : boolean;
  signal type_cast_1131_inst_req_0 : boolean;
  signal type_cast_915_inst_req_0 : boolean;
  signal ptr_deref_1013_store_0_ack_1 : boolean;
  signal type_cast_624_inst_req_0 : boolean;
  signal type_cast_624_inst_ack_0 : boolean;
  signal addr_of_877_final_reg_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_570_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_595_inst_req_0 : boolean;
  signal addr_of_877_final_reg_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_570_inst_ack_0 : boolean;
  signal if_stmt_1539_branch_ack_0 : boolean;
  signal type_cast_933_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_582_inst_ack_1 : boolean;
  signal type_cast_969_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_595_inst_ack_1 : boolean;
  signal type_cast_599_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_557_inst_ack_0 : boolean;
  signal type_cast_933_inst_ack_0 : boolean;
  signal type_cast_561_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_595_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_570_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_557_inst_ack_1 : boolean;
  signal if_stmt_1153_branch_ack_1 : boolean;
  signal type_cast_561_inst_req_1 : boolean;
  signal type_cast_599_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_557_inst_req_1 : boolean;
  signal if_stmt_1027_branch_req_0 : boolean;
  signal type_cast_599_inst_req_1 : boolean;
  signal type_cast_969_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_620_inst_req_0 : boolean;
  signal type_cast_915_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_620_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_557_inst_req_0 : boolean;
  signal type_cast_884_inst_ack_0 : boolean;
  signal array_obj_ref_876_index_offset_ack_0 : boolean;
  signal array_obj_ref_876_index_offset_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_607_inst_req_0 : boolean;
  signal type_cast_969_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_607_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1001_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_607_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_607_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_582_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_582_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_582_inst_req_0 : boolean;
  signal type_cast_611_inst_req_1 : boolean;
  signal type_cast_611_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_1723_inst_ack_0 : boolean;
  signal type_cast_1131_inst_ack_0 : boolean;
  signal type_cast_574_inst_req_1 : boolean;
  signal type_cast_915_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_595_inst_ack_0 : boolean;
  signal type_cast_561_inst_req_0 : boolean;
  signal type_cast_915_inst_ack_1 : boolean;
  signal type_cast_574_inst_ack_0 : boolean;
  signal type_cast_574_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1001_inst_ack_1 : boolean;
  signal type_cast_1131_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1001_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_929_inst_ack_1 : boolean;
  signal type_cast_1131_inst_req_1 : boolean;
  signal if_stmt_1153_branch_req_0 : boolean;
  signal type_cast_586_inst_req_0 : boolean;
  signal type_cast_586_inst_ack_1 : boolean;
  signal type_cast_611_inst_ack_0 : boolean;
  signal ptr_deref_1013_store_0_ack_0 : boolean;
  signal if_stmt_1078_branch_ack_1 : boolean;
  signal type_cast_611_inst_req_0 : boolean;
  signal type_cast_884_inst_ack_1 : boolean;
  signal type_cast_624_inst_req_1 : boolean;
  signal type_cast_624_inst_ack_1 : boolean;
  signal if_stmt_1488_branch_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_632_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_965_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_632_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_632_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_965_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_632_inst_ack_1 : boolean;
  signal ptr_deref_1013_store_0_req_1 : boolean;
  signal type_cast_636_inst_req_0 : boolean;
  signal type_cast_636_inst_ack_0 : boolean;
  signal if_stmt_1078_branch_req_0 : boolean;
  signal type_cast_636_inst_req_1 : boolean;
  signal type_cast_636_inst_ack_1 : boolean;
  signal type_cast_1146_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_645_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_965_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_645_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_645_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_965_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_645_inst_ack_1 : boolean;
  signal if_stmt_1153_branch_ack_0 : boolean;
  signal type_cast_987_inst_ack_1 : boolean;
  signal type_cast_987_inst_req_1 : boolean;
  signal type_cast_649_inst_req_0 : boolean;
  signal type_cast_649_inst_ack_0 : boolean;
  signal type_cast_649_inst_req_1 : boolean;
  signal type_cast_649_inst_ack_1 : boolean;
  signal type_cast_1146_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_657_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_657_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_657_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_657_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1127_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_911_inst_ack_1 : boolean;
  signal type_cast_661_inst_req_0 : boolean;
  signal type_cast_661_inst_ack_0 : boolean;
  signal type_cast_661_inst_req_1 : boolean;
  signal type_cast_951_inst_ack_1 : boolean;
  signal type_cast_661_inst_ack_1 : boolean;
  signal type_cast_1691_inst_ack_1 : boolean;
  signal type_cast_987_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_670_inst_req_0 : boolean;
  signal type_cast_951_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_670_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_670_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_670_inst_ack_1 : boolean;
  signal type_cast_1774_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1127_inst_req_1 : boolean;
  signal type_cast_987_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_911_inst_req_1 : boolean;
  signal type_cast_674_inst_req_0 : boolean;
  signal type_cast_674_inst_ack_0 : boolean;
  signal type_cast_674_inst_req_1 : boolean;
  signal type_cast_951_inst_ack_0 : boolean;
  signal type_cast_674_inst_ack_1 : boolean;
  signal type_cast_1146_inst_ack_0 : boolean;
  signal type_cast_1146_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_682_inst_req_0 : boolean;
  signal type_cast_951_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_682_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_880_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_682_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_682_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1127_inst_ack_0 : boolean;
  signal type_cast_686_inst_req_0 : boolean;
  signal type_cast_686_inst_ack_0 : boolean;
  signal type_cast_686_inst_req_1 : boolean;
  signal type_cast_686_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_695_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_695_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_880_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_695_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_695_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1127_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_911_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_911_inst_req_0 : boolean;
  signal type_cast_699_inst_req_0 : boolean;
  signal type_cast_699_inst_ack_0 : boolean;
  signal type_cast_699_inst_req_1 : boolean;
  signal type_cast_699_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_707_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_947_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_707_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_880_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_707_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_947_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_707_inst_ack_1 : boolean;
  signal type_cast_897_inst_ack_1 : boolean;
  signal type_cast_897_inst_req_1 : boolean;
  signal if_stmt_1027_branch_ack_0 : boolean;
  signal type_cast_711_inst_req_0 : boolean;
  signal type_cast_711_inst_ack_0 : boolean;
  signal type_cast_711_inst_req_1 : boolean;
  signal type_cast_711_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_880_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_983_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_983_inst_req_1 : boolean;
  signal type_cast_1005_inst_ack_1 : boolean;
  signal type_cast_1005_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_720_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_947_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_720_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_720_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_947_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_720_inst_ack_1 : boolean;
  signal type_cast_897_inst_ack_0 : boolean;
  signal type_cast_897_inst_req_0 : boolean;
  signal type_cast_724_inst_req_0 : boolean;
  signal type_cast_724_inst_ack_0 : boolean;
  signal if_stmt_1027_branch_ack_1 : boolean;
  signal type_cast_724_inst_req_1 : boolean;
  signal type_cast_724_inst_ack_1 : boolean;
  signal type_cast_1005_inst_ack_0 : boolean;
  signal type_cast_1005_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_732_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_732_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_732_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_732_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_893_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_893_inst_req_1 : boolean;
  signal type_cast_736_inst_req_0 : boolean;
  signal type_cast_736_inst_ack_0 : boolean;
  signal type_cast_736_inst_req_1 : boolean;
  signal type_cast_736_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_983_inst_ack_0 : boolean;
  signal addr_of_877_final_reg_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_983_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_745_inst_req_0 : boolean;
  signal type_cast_933_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_745_inst_ack_0 : boolean;
  signal addr_of_877_final_reg_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_745_inst_req_1 : boolean;
  signal type_cast_933_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_745_inst_ack_1 : boolean;
  signal type_cast_749_inst_req_0 : boolean;
  signal type_cast_749_inst_ack_0 : boolean;
  signal type_cast_749_inst_req_1 : boolean;
  signal type_cast_749_inst_ack_1 : boolean;
  signal type_cast_758_inst_req_0 : boolean;
  signal call_stmt_1668_call_req_0 : boolean;
  signal type_cast_758_inst_ack_0 : boolean;
  signal if_stmt_1488_branch_ack_1 : boolean;
  signal if_stmt_1753_branch_req_0 : boolean;
  signal type_cast_758_inst_req_1 : boolean;
  signal type_cast_758_inst_ack_1 : boolean;
  signal if_stmt_1488_branch_ack_0 : boolean;
  signal type_cast_762_inst_req_0 : boolean;
  signal call_stmt_1668_call_ack_0 : boolean;
  signal type_cast_762_inst_ack_0 : boolean;
  signal type_cast_762_inst_req_1 : boolean;
  signal type_cast_762_inst_ack_1 : boolean;
  signal type_cast_778_inst_req_0 : boolean;
  signal type_cast_778_inst_ack_0 : boolean;
  signal type_cast_778_inst_req_1 : boolean;
  signal type_cast_778_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_1726_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1592_inst_req_0 : boolean;
  signal WPIPE_num_out_pipe_1723_inst_req_1 : boolean;
  signal WPIPE_num_out_pipe_1723_inst_ack_1 : boolean;
  signal if_stmt_1753_branch_ack_1 : boolean;
  signal if_stmt_786_branch_req_0 : boolean;
  signal array_obj_ref_1657_index_offset_req_0 : boolean;
  signal if_stmt_786_branch_ack_1 : boolean;
  signal if_stmt_786_branch_ack_0 : boolean;
  signal type_cast_806_inst_req_0 : boolean;
  signal type_cast_806_inst_ack_0 : boolean;
  signal type_cast_806_inst_req_1 : boolean;
  signal type_cast_806_inst_ack_1 : boolean;
  signal type_cast_822_inst_req_0 : boolean;
  signal type_cast_822_inst_ack_0 : boolean;
  signal type_cast_822_inst_req_1 : boolean;
  signal type_cast_822_inst_ack_1 : boolean;
  signal type_cast_831_inst_req_0 : boolean;
  signal type_cast_831_inst_ack_0 : boolean;
  signal type_cast_831_inst_req_1 : boolean;
  signal type_cast_831_inst_ack_1 : boolean;
  signal type_cast_841_inst_req_0 : boolean;
  signal type_cast_841_inst_ack_0 : boolean;
  signal type_cast_841_inst_req_1 : boolean;
  signal type_cast_841_inst_ack_1 : boolean;
  signal array_obj_ref_1192_index_offset_ack_0 : boolean;
  signal array_obj_ref_1192_index_offset_req_1 : boolean;
  signal array_obj_ref_1192_index_offset_ack_1 : boolean;
  signal WPIPE_num_out_pipe_1726_inst_req_0 : boolean;
  signal type_cast_1774_inst_ack_1 : boolean;
  signal RPIPE_input_done_pipe_1766_inst_req_0 : boolean;
  signal addr_of_1193_final_reg_req_0 : boolean;
  signal addr_of_1193_final_reg_ack_0 : boolean;
  signal addr_of_1193_final_reg_req_1 : boolean;
  signal addr_of_1193_final_reg_ack_1 : boolean;
  signal type_cast_1774_inst_req_0 : boolean;
  signal call_stmt_1770_call_ack_1 : boolean;
  signal call_stmt_1770_call_req_1 : boolean;
  signal type_cast_1691_inst_req_1 : boolean;
  signal type_cast_1691_inst_ack_0 : boolean;
  signal type_cast_1691_inst_req_0 : boolean;
  signal ptr_deref_1661_store_0_ack_1 : boolean;
  signal ptr_deref_1661_store_0_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1592_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_1723_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1592_inst_req_1 : boolean;
  signal ptr_deref_1196_store_0_req_0 : boolean;
  signal ptr_deref_1196_store_0_ack_0 : boolean;
  signal ptr_deref_1196_store_0_req_1 : boolean;
  signal ptr_deref_1196_store_0_ack_1 : boolean;
  signal type_cast_1203_inst_req_0 : boolean;
  signal type_cast_1203_inst_ack_0 : boolean;
  signal type_cast_1203_inst_req_1 : boolean;
  signal type_cast_1203_inst_ack_1 : boolean;
  signal call_stmt_1770_call_ack_0 : boolean;
  signal call_stmt_1770_call_req_0 : boolean;
  signal type_cast_1207_inst_req_0 : boolean;
  signal type_cast_1207_inst_ack_0 : boolean;
  signal type_cast_1207_inst_req_1 : boolean;
  signal type_cast_1207_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1674_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1674_inst_req_1 : boolean;
  signal if_stmt_1753_branch_ack_0 : boolean;
  signal type_cast_1211_inst_req_0 : boolean;
  signal ptr_deref_1661_store_0_ack_0 : boolean;
  signal type_cast_1211_inst_ack_0 : boolean;
  signal call_stmt_1741_call_ack_1 : boolean;
  signal type_cast_1211_inst_req_1 : boolean;
  signal ptr_deref_1661_store_0_req_0 : boolean;
  signal type_cast_1211_inst_ack_1 : boolean;
  signal type_cast_1783_inst_req_0 : boolean;
  signal type_cast_1783_inst_ack_0 : boolean;
  signal call_stmt_1741_call_req_1 : boolean;
  signal type_cast_1774_inst_req_1 : boolean;
  signal if_stmt_1539_branch_ack_1 : boolean;
  signal if_stmt_1249_branch_req_0 : boolean;
  signal array_obj_ref_1657_index_offset_ack_1 : boolean;
  signal if_stmt_1249_branch_ack_1 : boolean;
  signal array_obj_ref_1657_index_offset_req_1 : boolean;
  signal if_stmt_1539_branch_req_0 : boolean;
  signal if_stmt_1249_branch_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1674_inst_ack_0 : boolean;
  signal type_cast_1270_inst_req_0 : boolean;
  signal type_cast_1270_inst_ack_0 : boolean;
  signal call_stmt_1741_call_ack_0 : boolean;
  signal call_stmt_1741_call_req_0 : boolean;
  signal type_cast_1270_inst_req_1 : boolean;
  signal type_cast_1270_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1674_inst_req_0 : boolean;
  signal type_cast_1279_inst_req_0 : boolean;
  signal type_cast_1279_inst_ack_0 : boolean;
  signal type_cast_1279_inst_req_1 : boolean;
  signal type_cast_1279_inst_ack_1 : boolean;
  signal type_cast_1288_inst_req_0 : boolean;
  signal type_cast_1288_inst_ack_0 : boolean;
  signal type_cast_1288_inst_req_1 : boolean;
  signal type_cast_1288_inst_ack_1 : boolean;
  signal RPIPE_input_done_pipe_1766_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1670_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1670_inst_req_1 : boolean;
  signal call_stmt_1737_call_ack_1 : boolean;
  signal type_cast_1297_inst_req_0 : boolean;
  signal type_cast_1297_inst_ack_0 : boolean;
  signal call_stmt_1737_call_req_1 : boolean;
  signal type_cast_1297_inst_req_1 : boolean;
  signal type_cast_1297_inst_ack_1 : boolean;
  signal RPIPE_input_done_pipe_1766_inst_req_1 : boolean;
  signal type_cast_1302_inst_req_0 : boolean;
  signal type_cast_1302_inst_ack_0 : boolean;
  signal call_stmt_1737_call_ack_0 : boolean;
  signal type_cast_1302_inst_req_1 : boolean;
  signal type_cast_1302_inst_ack_1 : boolean;
  signal RPIPE_input_done_pipe_1766_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1670_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1670_inst_req_0 : boolean;
  signal array_obj_ref_1657_index_offset_ack_0 : boolean;
  signal call_stmt_1737_call_req_0 : boolean;
  signal if_stmt_1618_branch_ack_0 : boolean;
  signal array_obj_ref_1337_index_offset_req_0 : boolean;
  signal array_obj_ref_1337_index_offset_ack_0 : boolean;
  signal array_obj_ref_1337_index_offset_req_1 : boolean;
  signal array_obj_ref_1337_index_offset_ack_1 : boolean;
  signal type_cast_1763_inst_ack_1 : boolean;
  signal addr_of_1338_final_reg_req_0 : boolean;
  signal addr_of_1338_final_reg_ack_0 : boolean;
  signal addr_of_1338_final_reg_req_1 : boolean;
  signal addr_of_1338_final_reg_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1341_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1341_inst_ack_0 : boolean;
  signal type_cast_1554_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1341_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1341_inst_ack_1 : boolean;
  signal type_cast_1763_inst_req_1 : boolean;
  signal if_stmt_1618_branch_ack_1 : boolean;
  signal if_stmt_1618_branch_req_0 : boolean;
  signal type_cast_1345_inst_req_0 : boolean;
  signal type_cast_1345_inst_ack_0 : boolean;
  signal type_cast_1345_inst_req_1 : boolean;
  signal type_cast_1345_inst_ack_1 : boolean;
  signal type_cast_1554_inst_req_1 : boolean;
  signal type_cast_1701_inst_ack_1 : boolean;
  signal type_cast_1701_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1592_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1354_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1354_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1354_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1354_inst_ack_1 : boolean;
  signal type_cast_1763_inst_ack_0 : boolean;
  signal type_cast_1611_inst_ack_1 : boolean;
  signal type_cast_1611_inst_req_1 : boolean;
  signal type_cast_1358_inst_req_0 : boolean;
  signal type_cast_1358_inst_ack_0 : boolean;
  signal type_cast_1358_inst_req_1 : boolean;
  signal type_cast_1358_inst_ack_1 : boolean;
  signal type_cast_1554_inst_ack_0 : boolean;
  signal type_cast_1554_inst_req_0 : boolean;
  signal call_stmt_1668_call_ack_1 : boolean;
  signal type_cast_1701_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1372_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1372_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1372_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1372_inst_ack_1 : boolean;
  signal type_cast_1763_inst_req_0 : boolean;
  signal type_cast_1611_inst_ack_0 : boolean;
  signal type_cast_1611_inst_req_0 : boolean;
  signal type_cast_1376_inst_req_0 : boolean;
  signal type_cast_1376_inst_ack_0 : boolean;
  signal type_cast_1376_inst_req_1 : boolean;
  signal type_cast_1376_inst_ack_1 : boolean;
  signal call_stmt_1668_call_req_1 : boolean;
  signal type_cast_1701_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1390_inst_req_0 : boolean;
  signal addr_of_1658_final_reg_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1390_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1390_inst_req_1 : boolean;
  signal addr_of_1658_final_reg_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1390_inst_ack_1 : boolean;
  signal type_cast_1596_inst_ack_1 : boolean;
  signal type_cast_1596_inst_req_1 : boolean;
  signal WPIPE_num_out_pipe_1726_inst_ack_1 : boolean;
  signal type_cast_1394_inst_req_0 : boolean;
  signal type_cast_1394_inst_ack_0 : boolean;
  signal type_cast_1394_inst_req_1 : boolean;
  signal type_cast_1394_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1408_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1408_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1408_inst_req_1 : boolean;
  signal addr_of_1658_final_reg_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1408_inst_ack_1 : boolean;
  signal type_cast_1596_inst_ack_0 : boolean;
  signal type_cast_1596_inst_req_0 : boolean;
  signal WPIPE_num_out_pipe_1726_inst_req_1 : boolean;
  signal type_cast_1412_inst_req_0 : boolean;
  signal addr_of_1658_final_reg_req_0 : boolean;
  signal type_cast_1412_inst_ack_0 : boolean;
  signal type_cast_1412_inst_req_1 : boolean;
  signal type_cast_1412_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1426_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1426_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1426_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1426_inst_ack_1 : boolean;
  signal type_cast_1430_inst_req_0 : boolean;
  signal type_cast_1430_inst_ack_0 : boolean;
  signal type_cast_1430_inst_req_1 : boolean;
  signal type_cast_1430_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1444_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1444_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1444_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1444_inst_ack_1 : boolean;
  signal type_cast_1448_inst_req_0 : boolean;
  signal type_cast_1448_inst_ack_0 : boolean;
  signal type_cast_1448_inst_req_1 : boolean;
  signal type_cast_1448_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1462_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1462_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1462_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1462_inst_ack_1 : boolean;
  signal type_cast_1466_inst_req_0 : boolean;
  signal type_cast_1466_inst_ack_0 : boolean;
  signal type_cast_1466_inst_req_1 : boolean;
  signal type_cast_1466_inst_ack_1 : boolean;
  signal ptr_deref_1474_store_0_req_0 : boolean;
  signal ptr_deref_1474_store_0_ack_0 : boolean;
  signal ptr_deref_1474_store_0_req_1 : boolean;
  signal ptr_deref_1474_store_0_ack_1 : boolean;
  signal type_cast_1783_inst_req_1 : boolean;
  signal type_cast_1783_inst_ack_1 : boolean;
  signal type_cast_1793_inst_req_0 : boolean;
  signal type_cast_1793_inst_ack_0 : boolean;
  signal type_cast_1793_inst_req_1 : boolean;
  signal type_cast_1793_inst_ack_1 : boolean;
  signal type_cast_1803_inst_req_0 : boolean;
  signal type_cast_1803_inst_ack_0 : boolean;
  signal type_cast_1803_inst_req_1 : boolean;
  signal type_cast_1803_inst_ack_1 : boolean;
  signal type_cast_1813_inst_req_0 : boolean;
  signal type_cast_1813_inst_ack_0 : boolean;
  signal type_cast_1813_inst_req_1 : boolean;
  signal type_cast_1813_inst_ack_1 : boolean;
  signal phi_stmt_1710_ack_0 : boolean;
  signal type_cast_1823_inst_req_0 : boolean;
  signal type_cast_1823_inst_ack_0 : boolean;
  signal type_cast_1823_inst_req_1 : boolean;
  signal type_cast_1823_inst_ack_1 : boolean;
  signal type_cast_1833_inst_req_0 : boolean;
  signal type_cast_1833_inst_ack_0 : boolean;
  signal type_cast_1833_inst_req_1 : boolean;
  signal type_cast_1833_inst_ack_1 : boolean;
  signal type_cast_1843_inst_req_0 : boolean;
  signal type_cast_1843_inst_ack_0 : boolean;
  signal type_cast_1843_inst_req_1 : boolean;
  signal type_cast_1843_inst_ack_1 : boolean;
  signal type_cast_1853_inst_req_0 : boolean;
  signal type_cast_1853_inst_ack_0 : boolean;
  signal type_cast_1853_inst_req_1 : boolean;
  signal type_cast_1853_inst_ack_1 : boolean;
  signal phi_stmt_1710_req_0 : boolean;
  signal type_cast_1713_inst_ack_1 : boolean;
  signal type_cast_1713_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1855_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1855_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1855_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1855_inst_ack_1 : boolean;
  signal phi_stmt_1564_req_1 : boolean;
  signal type_cast_1570_inst_ack_1 : boolean;
  signal type_cast_1570_inst_req_1 : boolean;
  signal type_cast_1570_inst_ack_0 : boolean;
  signal type_cast_1570_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1858_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1858_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1858_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1858_inst_ack_1 : boolean;
  signal type_cast_1713_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1861_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1861_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1861_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1861_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1864_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1864_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1864_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1864_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1867_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1867_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1867_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1867_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1870_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1870_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1870_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1870_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1873_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1873_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1873_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1873_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1876_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1876_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1876_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1876_inst_ack_1 : boolean;
  signal type_cast_1713_inst_req_0 : boolean;
  signal phi_stmt_864_req_0 : boolean;
  signal type_cast_870_inst_req_0 : boolean;
  signal type_cast_870_inst_ack_0 : boolean;
  signal type_cast_870_inst_req_1 : boolean;
  signal type_cast_870_inst_ack_1 : boolean;
  signal phi_stmt_864_req_1 : boolean;
  signal phi_stmt_864_ack_0 : boolean;
  signal phi_stmt_1625_ack_0 : boolean;
  signal phi_stmt_1058_req_1 : boolean;
  signal type_cast_1061_inst_req_0 : boolean;
  signal type_cast_1061_inst_ack_0 : boolean;
  signal type_cast_1061_inst_req_1 : boolean;
  signal type_cast_1061_inst_ack_1 : boolean;
  signal phi_stmt_1058_req_0 : boolean;
  signal phi_stmt_1571_ack_0 : boolean;
  signal phi_stmt_1058_ack_0 : boolean;
  signal phi_stmt_1564_ack_0 : boolean;
  signal phi_stmt_1099_req_0 : boolean;
  signal phi_stmt_1106_req_0 : boolean;
  signal type_cast_1105_inst_req_0 : boolean;
  signal type_cast_1105_inst_ack_0 : boolean;
  signal type_cast_1105_inst_req_1 : boolean;
  signal type_cast_1105_inst_ack_1 : boolean;
  signal phi_stmt_1099_req_1 : boolean;
  signal phi_stmt_1571_req_1 : boolean;
  signal phi_stmt_1625_req_0 : boolean;
  signal type_cast_1112_inst_req_0 : boolean;
  signal type_cast_1112_inst_ack_0 : boolean;
  signal type_cast_1112_inst_req_1 : boolean;
  signal type_cast_1112_inst_ack_1 : boolean;
  signal phi_stmt_1106_req_1 : boolean;
  signal phi_stmt_1099_ack_0 : boolean;
  signal phi_stmt_1106_ack_0 : boolean;
  signal type_cast_1577_inst_ack_1 : boolean;
  signal type_cast_1628_inst_ack_1 : boolean;
  signal phi_stmt_1710_req_1 : boolean;
  signal type_cast_1628_inst_req_1 : boolean;
  signal type_cast_1163_inst_req_0 : boolean;
  signal type_cast_1163_inst_ack_0 : boolean;
  signal type_cast_1163_inst_req_1 : boolean;
  signal type_cast_1163_inst_ack_1 : boolean;
  signal phi_stmt_1160_req_0 : boolean;
  signal phi_stmt_1571_req_0 : boolean;
  signal phi_stmt_1160_ack_0 : boolean;
  signal type_cast_1577_inst_req_1 : boolean;
  signal phi_stmt_1325_req_0 : boolean;
  signal type_cast_1331_inst_req_0 : boolean;
  signal type_cast_1331_inst_ack_0 : boolean;
  signal type_cast_1331_inst_req_1 : boolean;
  signal type_cast_1331_inst_ack_1 : boolean;
  signal phi_stmt_1325_req_1 : boolean;
  signal phi_stmt_1325_ack_0 : boolean;
  signal type_cast_1577_inst_ack_0 : boolean;
  signal type_cast_1577_inst_req_0 : boolean;
  signal type_cast_1628_inst_ack_0 : boolean;
  signal type_cast_1522_inst_req_0 : boolean;
  signal type_cast_1522_inst_ack_0 : boolean;
  signal type_cast_1522_inst_req_1 : boolean;
  signal type_cast_1522_inst_ack_1 : boolean;
  signal phi_stmt_1519_req_0 : boolean;
  signal phi_stmt_1519_req_1 : boolean;
  signal phi_stmt_1519_ack_0 : boolean;
  signal type_cast_1628_inst_req_0 : boolean;
  signal phi_stmt_1564_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolution3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolution3D_CP_1767_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolution3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_1767_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolution3D_CP_1767_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_1767_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolution3D_CP_1767: Block -- control-path 
    signal convolution3D_CP_1767_elements: BooleanArray(366 downto 0);
    -- 
  begin -- 
    convolution3D_CP_1767_elements(0) <= convolution3D_CP_1767_start;
    convolution3D_CP_1767_symbol <= convolution3D_CP_1767_elements(298);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	64 
    -- CP-element group 0: 	67 
    -- CP-element group 0: 	70 
    -- CP-element group 0: 	73 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0:  members (65) 
      -- CP-element group 0: 	 branch_block_stmt_554/branch_block_stmt_554__entry__
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_599_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_557_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_586_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_624_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_624_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_611_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_557_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_554/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_561_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_599_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785__entry__
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_561_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_557_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_611_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_611_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_586_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_574_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_574_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_586_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_574_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_599_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_561_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_624_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_636_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_636_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_636_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_649_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_649_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_649_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_661_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_661_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_661_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_674_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_674_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_674_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_686_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_686_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_686_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_699_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_699_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_699_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_711_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_711_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_711_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_724_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_724_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_724_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_736_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_736_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_736_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_749_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_749_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_749_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_758_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_758_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_758_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_762_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_762_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_762_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_778_update_start_
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_778_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_778_Update/cr
      -- 
    cr_1958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_586_inst_req_1); -- 
    cr_1902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_561_inst_req_1); -- 
    cr_1986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_599_inst_req_1); -- 
    rr_1883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => RPIPE_maxpool_input_pipe_557_inst_req_0); -- 
    cr_2014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_611_inst_req_1); -- 
    cr_1930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_574_inst_req_1); -- 
    cr_2042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_624_inst_req_1); -- 
    cr_2070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_636_inst_req_1); -- 
    cr_2098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_649_inst_req_1); -- 
    cr_2126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_661_inst_req_1); -- 
    cr_2154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_674_inst_req_1); -- 
    cr_2182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_686_inst_req_1); -- 
    cr_2210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_699_inst_req_1); -- 
    cr_2238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_711_inst_req_1); -- 
    cr_2266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_724_inst_req_1); -- 
    cr_2294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_736_inst_req_1); -- 
    cr_2322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_749_inst_req_1); -- 
    cr_2336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_758_inst_req_1); -- 
    cr_2350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_762_inst_req_1); -- 
    cr_2364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(0), ack => type_cast_778_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_557_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_557_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_557_update_start_
      -- CP-element group 1: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_557_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_557_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_557_Update/cr
      -- 
    ra_1884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_557_inst_ack_0, ack => convolution3D_CP_1767_elements(1)); -- 
    cr_1888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(1), ack => RPIPE_maxpool_input_pipe_557_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_557_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_561_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_570_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_570_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_557_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_557_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_570_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_561_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_561_Sample/$entry
      -- 
    ca_1889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_557_inst_ack_1, ack => convolution3D_CP_1767_elements(2)); -- 
    rr_1897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(2), ack => type_cast_561_inst_req_0); -- 
    rr_1911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(2), ack => RPIPE_maxpool_input_pipe_570_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_561_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_561_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_561_Sample/$exit
      -- 
    ra_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_561_inst_ack_0, ack => convolution3D_CP_1767_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	71 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_561_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_561_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_561_update_completed_
      -- 
    ca_1903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_561_inst_ack_1, ack => convolution3D_CP_1767_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_570_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_570_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_570_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_570_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_570_update_start_
      -- CP-element group 5: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_570_sample_completed_
      -- 
    ra_1912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_570_inst_ack_0, ack => convolution3D_CP_1767_elements(5)); -- 
    cr_1916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(5), ack => RPIPE_maxpool_input_pipe_570_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_570_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_570_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_570_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_582_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_582_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_582_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_574_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_574_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_574_sample_start_
      -- 
    ca_1917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_570_inst_ack_1, ack => convolution3D_CP_1767_elements(6)); -- 
    rr_1925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(6), ack => type_cast_574_inst_req_0); -- 
    rr_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(6), ack => RPIPE_maxpool_input_pipe_582_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_574_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_574_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_574_sample_completed_
      -- 
    ra_1926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_574_inst_ack_0, ack => convolution3D_CP_1767_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	71 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_574_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_574_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_574_update_completed_
      -- 
    ca_1931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_574_inst_ack_1, ack => convolution3D_CP_1767_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_582_update_start_
      -- CP-element group 9: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_582_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_582_Update/cr
      -- CP-element group 9: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_582_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_582_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_582_Sample/$exit
      -- 
    ra_1940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_582_inst_ack_0, ack => convolution3D_CP_1767_elements(9)); -- 
    cr_1944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(9), ack => RPIPE_maxpool_input_pipe_582_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_595_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_595_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_582_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_582_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_582_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_586_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_595_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_586_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_586_Sample/rr
      -- 
    ca_1945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_582_inst_ack_1, ack => convolution3D_CP_1767_elements(10)); -- 
    rr_1953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(10), ack => type_cast_586_inst_req_0); -- 
    rr_1967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(10), ack => RPIPE_maxpool_input_pipe_595_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_586_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_586_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_586_Sample/$exit
      -- 
    ra_1954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_586_inst_ack_0, ack => convolution3D_CP_1767_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	65 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_586_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_586_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_586_Update/ca
      -- 
    ca_1959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_586_inst_ack_1, ack => convolution3D_CP_1767_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_595_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_595_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_595_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_595_update_start_
      -- CP-element group 13: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_595_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_595_sample_completed_
      -- 
    ra_1968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_595_inst_ack_0, ack => convolution3D_CP_1767_elements(13)); -- 
    cr_1972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(13), ack => RPIPE_maxpool_input_pipe_595_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_595_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_599_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_599_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_595_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_607_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_595_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_599_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_607_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_607_Sample/$entry
      -- 
    ca_1973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_595_inst_ack_1, ack => convolution3D_CP_1767_elements(14)); -- 
    rr_1981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(14), ack => type_cast_599_inst_req_0); -- 
    rr_1995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(14), ack => RPIPE_maxpool_input_pipe_607_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_599_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_599_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_599_Sample/$exit
      -- 
    ra_1982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_599_inst_ack_0, ack => convolution3D_CP_1767_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	65 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_599_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_599_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_599_update_completed_
      -- 
    ca_1987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_599_inst_ack_1, ack => convolution3D_CP_1767_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_607_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_607_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_607_Update/cr
      -- CP-element group 17: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_607_update_start_
      -- CP-element group 17: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_607_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_607_Sample/$exit
      -- 
    ra_1996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_607_inst_ack_0, ack => convolution3D_CP_1767_elements(17)); -- 
    cr_2000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(17), ack => RPIPE_maxpool_input_pipe_607_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_620_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_620_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_620_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_607_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_611_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_607_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_611_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_607_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_611_Sample/rr
      -- 
    ca_2001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_607_inst_ack_1, ack => convolution3D_CP_1767_elements(18)); -- 
    rr_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(18), ack => type_cast_611_inst_req_0); -- 
    rr_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(18), ack => RPIPE_maxpool_input_pipe_620_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_611_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_611_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_611_Sample/$exit
      -- 
    ra_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_611_inst_ack_0, ack => convolution3D_CP_1767_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	68 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_611_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_611_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_611_Update/ca
      -- 
    ca_2015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_611_inst_ack_1, ack => convolution3D_CP_1767_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_620_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_620_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_620_update_start_
      -- CP-element group 21: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_620_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_620_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_620_Sample/ra
      -- 
    ra_2024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_620_inst_ack_0, ack => convolution3D_CP_1767_elements(21)); -- 
    cr_2028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(21), ack => RPIPE_maxpool_input_pipe_620_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	25 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_620_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_620_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_620_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_624_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_624_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_624_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_632_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_632_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_632_Sample/rr
      -- 
    ca_2029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_620_inst_ack_1, ack => convolution3D_CP_1767_elements(22)); -- 
    rr_2037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(22), ack => type_cast_624_inst_req_0); -- 
    rr_2051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(22), ack => RPIPE_maxpool_input_pipe_632_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_624_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_624_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_624_Sample/ra
      -- 
    ra_2038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_624_inst_ack_0, ack => convolution3D_CP_1767_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	68 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_624_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_624_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_624_Update/ca
      -- 
    ca_2043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_624_inst_ack_1, ack => convolution3D_CP_1767_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_632_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_632_update_start_
      -- CP-element group 25: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_632_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_632_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_632_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_632_Update/cr
      -- 
    ra_2052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_632_inst_ack_0, ack => convolution3D_CP_1767_elements(25)); -- 
    cr_2056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(25), ack => RPIPE_maxpool_input_pipe_632_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_632_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_632_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_632_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_636_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_636_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_636_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_645_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_645_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_645_Sample/rr
      -- 
    ca_2057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_632_inst_ack_1, ack => convolution3D_CP_1767_elements(26)); -- 
    rr_2065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(26), ack => type_cast_636_inst_req_0); -- 
    rr_2079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(26), ack => RPIPE_maxpool_input_pipe_645_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_636_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_636_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_636_Sample/ra
      -- 
    ra_2066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_636_inst_ack_0, ack => convolution3D_CP_1767_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	74 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_636_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_636_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_636_Update/ca
      -- 
    ca_2071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_636_inst_ack_1, ack => convolution3D_CP_1767_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_645_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_645_update_start_
      -- CP-element group 29: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_645_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_645_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_645_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_645_Update/cr
      -- 
    ra_2080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_645_inst_ack_0, ack => convolution3D_CP_1767_elements(29)); -- 
    cr_2084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(29), ack => RPIPE_maxpool_input_pipe_645_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_645_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_645_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_645_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_649_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_649_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_649_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_657_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_657_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_657_Sample/rr
      -- 
    ca_2085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_645_inst_ack_1, ack => convolution3D_CP_1767_elements(30)); -- 
    rr_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(30), ack => type_cast_649_inst_req_0); -- 
    rr_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(30), ack => RPIPE_maxpool_input_pipe_657_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_649_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_649_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_649_Sample/ra
      -- 
    ra_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_649_inst_ack_0, ack => convolution3D_CP_1767_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	74 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_649_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_649_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_649_Update/ca
      -- 
    ca_2099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_649_inst_ack_1, ack => convolution3D_CP_1767_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_657_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_657_update_start_
      -- CP-element group 33: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_657_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_657_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_657_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_657_Update/cr
      -- 
    ra_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_657_inst_ack_0, ack => convolution3D_CP_1767_elements(33)); -- 
    cr_2112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(33), ack => RPIPE_maxpool_input_pipe_657_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_657_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_657_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_657_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_661_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_661_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_661_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_670_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_670_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_670_Sample/rr
      -- 
    ca_2113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_657_inst_ack_1, ack => convolution3D_CP_1767_elements(34)); -- 
    rr_2121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(34), ack => type_cast_661_inst_req_0); -- 
    rr_2135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(34), ack => RPIPE_maxpool_input_pipe_670_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_661_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_661_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_661_Sample/ra
      -- 
    ra_2122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_661_inst_ack_0, ack => convolution3D_CP_1767_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	74 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_661_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_661_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_661_Update/ca
      -- 
    ca_2127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_661_inst_ack_1, ack => convolution3D_CP_1767_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_670_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_670_update_start_
      -- CP-element group 37: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_670_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_670_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_670_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_670_Update/cr
      -- 
    ra_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_670_inst_ack_0, ack => convolution3D_CP_1767_elements(37)); -- 
    cr_2140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(37), ack => RPIPE_maxpool_input_pipe_670_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	41 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_670_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_670_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_670_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_674_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_674_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_674_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_682_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_682_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_682_Sample/rr
      -- 
    ca_2141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_670_inst_ack_1, ack => convolution3D_CP_1767_elements(38)); -- 
    rr_2163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(38), ack => RPIPE_maxpool_input_pipe_682_inst_req_0); -- 
    rr_2149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(38), ack => type_cast_674_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_674_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_674_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_674_Sample/ra
      -- 
    ra_2150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_674_inst_ack_0, ack => convolution3D_CP_1767_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	74 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_674_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_674_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_674_Update/ca
      -- 
    ca_2155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_674_inst_ack_1, ack => convolution3D_CP_1767_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_682_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_682_update_start_
      -- CP-element group 41: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_682_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_682_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_682_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_682_Update/cr
      -- 
    ra_2164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_682_inst_ack_0, ack => convolution3D_CP_1767_elements(41)); -- 
    cr_2168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(41), ack => RPIPE_maxpool_input_pipe_682_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_682_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_682_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_682_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_686_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_686_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_686_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_695_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_695_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_695_Sample/rr
      -- 
    ca_2169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_682_inst_ack_1, ack => convolution3D_CP_1767_elements(42)); -- 
    rr_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(42), ack => type_cast_686_inst_req_0); -- 
    rr_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(42), ack => RPIPE_maxpool_input_pipe_695_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_686_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_686_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_686_Sample/ra
      -- 
    ra_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_686_inst_ack_0, ack => convolution3D_CP_1767_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	74 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_686_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_686_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_686_Update/ca
      -- 
    ca_2183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_686_inst_ack_1, ack => convolution3D_CP_1767_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_695_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_695_update_start_
      -- CP-element group 45: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_695_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_695_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_695_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_695_Update/cr
      -- 
    ra_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_695_inst_ack_0, ack => convolution3D_CP_1767_elements(45)); -- 
    cr_2196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(45), ack => RPIPE_maxpool_input_pipe_695_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_695_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_695_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_695_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_699_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_699_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_699_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_707_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_707_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_707_Sample/rr
      -- 
    ca_2197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_695_inst_ack_1, ack => convolution3D_CP_1767_elements(46)); -- 
    rr_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(46), ack => type_cast_699_inst_req_0); -- 
    rr_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(46), ack => RPIPE_maxpool_input_pipe_707_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_699_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_699_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_699_Sample/ra
      -- 
    ra_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_699_inst_ack_0, ack => convolution3D_CP_1767_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	74 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_699_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_699_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_699_Update/ca
      -- 
    ca_2211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_699_inst_ack_1, ack => convolution3D_CP_1767_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_707_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_707_update_start_
      -- CP-element group 49: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_707_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_707_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_707_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_707_Update/cr
      -- 
    ra_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_707_inst_ack_0, ack => convolution3D_CP_1767_elements(49)); -- 
    cr_2224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(49), ack => RPIPE_maxpool_input_pipe_707_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_707_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_707_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_707_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_711_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_711_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_711_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_720_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_720_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_720_Sample/rr
      -- 
    ca_2225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_707_inst_ack_1, ack => convolution3D_CP_1767_elements(50)); -- 
    rr_2233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(50), ack => type_cast_711_inst_req_0); -- 
    rr_2247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(50), ack => RPIPE_maxpool_input_pipe_720_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_711_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_711_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_711_Sample/ra
      -- 
    ra_2234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_711_inst_ack_0, ack => convolution3D_CP_1767_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	74 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_711_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_711_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_711_Update/ca
      -- 
    ca_2239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_711_inst_ack_1, ack => convolution3D_CP_1767_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_720_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_720_update_start_
      -- CP-element group 53: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_720_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_720_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_720_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_720_Update/cr
      -- 
    ra_2248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_720_inst_ack_0, ack => convolution3D_CP_1767_elements(53)); -- 
    cr_2252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(53), ack => RPIPE_maxpool_input_pipe_720_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	57 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_720_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_720_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_720_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_724_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_724_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_724_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_732_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_732_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_732_Sample/rr
      -- 
    ca_2253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_720_inst_ack_1, ack => convolution3D_CP_1767_elements(54)); -- 
    rr_2261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(54), ack => type_cast_724_inst_req_0); -- 
    rr_2275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(54), ack => RPIPE_maxpool_input_pipe_732_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_724_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_724_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_724_Sample/ra
      -- 
    ra_2262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_724_inst_ack_0, ack => convolution3D_CP_1767_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	74 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_724_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_724_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_724_Update/ca
      -- 
    ca_2267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_724_inst_ack_1, ack => convolution3D_CP_1767_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_732_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_732_update_start_
      -- CP-element group 57: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_732_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_732_Sample/ra
      -- CP-element group 57: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_732_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_732_Update/cr
      -- 
    ra_2276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_732_inst_ack_0, ack => convolution3D_CP_1767_elements(57)); -- 
    cr_2280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(57), ack => RPIPE_maxpool_input_pipe_732_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	61 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_732_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_732_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_732_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_736_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_736_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_736_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_745_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_745_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_745_Sample/rr
      -- 
    ca_2281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_732_inst_ack_1, ack => convolution3D_CP_1767_elements(58)); -- 
    rr_2289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(58), ack => type_cast_736_inst_req_0); -- 
    rr_2303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(58), ack => RPIPE_maxpool_input_pipe_745_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_736_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_736_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_736_Sample/ra
      -- 
    ra_2290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_736_inst_ack_0, ack => convolution3D_CP_1767_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	74 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_736_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_736_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_736_Update/ca
      -- 
    ca_2295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_736_inst_ack_1, ack => convolution3D_CP_1767_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	58 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_745_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_745_update_start_
      -- CP-element group 61: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_745_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_745_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_745_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_745_Update/cr
      -- 
    ra_2304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_745_inst_ack_0, ack => convolution3D_CP_1767_elements(61)); -- 
    cr_2308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(61), ack => RPIPE_maxpool_input_pipe_745_inst_req_1); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_745_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_745_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/RPIPE_maxpool_input_pipe_745_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_749_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_749_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_749_Sample/rr
      -- 
    ca_2309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_745_inst_ack_1, ack => convolution3D_CP_1767_elements(62)); -- 
    rr_2317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(62), ack => type_cast_749_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_749_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_749_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_749_Sample/ra
      -- 
    ra_2318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_749_inst_ack_0, ack => convolution3D_CP_1767_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	0 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	74 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_749_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_749_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_749_Update/ca
      -- 
    ca_2323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_749_inst_ack_1, ack => convolution3D_CP_1767_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	12 
    -- CP-element group 65: 	16 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_758_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_758_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_758_Sample/rr
      -- 
    rr_2331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(65), ack => type_cast_758_inst_req_0); -- 
    convolution3D_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(12) & convolution3D_CP_1767_elements(16);
      gj_convolution3D_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_758_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_758_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_758_Sample/ra
      -- 
    ra_2332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_758_inst_ack_0, ack => convolution3D_CP_1767_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	0 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	71 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_758_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_758_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_758_Update/ca
      -- 
    ca_2337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_758_inst_ack_1, ack => convolution3D_CP_1767_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	20 
    -- CP-element group 68: 	24 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_762_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_762_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_762_Sample/rr
      -- 
    rr_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(68), ack => type_cast_762_inst_req_0); -- 
    convolution3D_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(20) & convolution3D_CP_1767_elements(24);
      gj_convolution3D_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_762_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_762_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_762_Sample/ra
      -- 
    ra_2346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_762_inst_ack_0, ack => convolution3D_CP_1767_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	0 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_762_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_762_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_762_Update/ca
      -- 
    ca_2351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_762_inst_ack_1, ack => convolution3D_CP_1767_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	67 
    -- CP-element group 71: 	70 
    -- CP-element group 71: 	4 
    -- CP-element group 71: 	8 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_778_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_778_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_778_Sample/rr
      -- 
    rr_2359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(71), ack => type_cast_778_inst_req_0); -- 
    convolution3D_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(67) & convolution3D_CP_1767_elements(70) & convolution3D_CP_1767_elements(4) & convolution3D_CP_1767_elements(8);
      gj_convolution3D_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_778_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_778_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_778_Sample/ra
      -- 
    ra_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_778_inst_ack_0, ack => convolution3D_CP_1767_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	0 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_778_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_778_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/type_cast_778_Update/ca
      -- 
    ca_2365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_778_inst_ack_1, ack => convolution3D_CP_1767_elements(73)); -- 
    -- CP-element group 74:  branch  join  transition  place  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	28 
    -- CP-element group 74: 	32 
    -- CP-element group 74: 	44 
    -- CP-element group 74: 	36 
    -- CP-element group 74: 	40 
    -- CP-element group 74: 	48 
    -- CP-element group 74: 	52 
    -- CP-element group 74: 	56 
    -- CP-element group 74: 	60 
    -- CP-element group 74: 	64 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (10) 
      -- CP-element group 74: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785/$exit
      -- CP-element group 74: 	 branch_block_stmt_554/if_stmt_786__entry__
      -- CP-element group 74: 	 branch_block_stmt_554/assign_stmt_558_to_assign_stmt_785__exit__
      -- CP-element group 74: 	 branch_block_stmt_554/if_stmt_786_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_554/if_stmt_786_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_554/if_stmt_786_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_554/if_stmt_786_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_554/R_cmp367_787_place
      -- CP-element group 74: 	 branch_block_stmt_554/if_stmt_786_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_554/if_stmt_786_else_link/$entry
      -- 
    branch_req_2373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(74), ack => if_stmt_786_branch_req_0); -- 
    convolution3D_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(28) & convolution3D_CP_1767_elements(32) & convolution3D_CP_1767_elements(44) & convolution3D_CP_1767_elements(36) & convolution3D_CP_1767_elements(40) & convolution3D_CP_1767_elements(48) & convolution3D_CP_1767_elements(52) & convolution3D_CP_1767_elements(56) & convolution3D_CP_1767_elements(60) & convolution3D_CP_1767_elements(64) & convolution3D_CP_1767_elements(73);
      gj_convolution3D_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: 	78 
    -- CP-element group 75: 	79 
    -- CP-element group 75: 	80 
    -- CP-element group 75: 	81 
    -- CP-element group 75: 	82 
    -- CP-element group 75: 	85 
    -- CP-element group 75:  members (33) 
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861__entry__
      -- CP-element group 75: 	 branch_block_stmt_554/merge_stmt_792__exit__
      -- CP-element group 75: 	 branch_block_stmt_554/if_stmt_786_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_554/if_stmt_786_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_554/entry_bbx_xnph369
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/$entry
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_806_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_806_update_start_
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_806_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_806_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_806_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_806_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_822_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_822_update_start_
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_822_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_822_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_822_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_822_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_831_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_831_update_start_
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_831_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_831_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_831_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_831_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_841_update_start_
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_841_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_841_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_554/entry_bbx_xnph369_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_554/entry_bbx_xnph369_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_554/merge_stmt_792_PhiReqMerge
      -- CP-element group 75: 	 branch_block_stmt_554/merge_stmt_792_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_554/merge_stmt_792_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_554/merge_stmt_792_PhiAck/dummy
      -- 
    if_choice_transition_2378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_786_branch_ack_1, ack => convolution3D_CP_1767_elements(75)); -- 
    rr_2395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(75), ack => type_cast_806_inst_req_0); -- 
    cr_2400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(75), ack => type_cast_806_inst_req_1); -- 
    rr_2409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(75), ack => type_cast_822_inst_req_0); -- 
    cr_2414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(75), ack => type_cast_822_inst_req_1); -- 
    rr_2423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(75), ack => type_cast_831_inst_req_0); -- 
    cr_2428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(75), ack => type_cast_831_inst_req_1); -- 
    cr_2442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(75), ack => type_cast_841_inst_req_1); -- 
    -- CP-element group 76:  transition  place  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	305 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_554/if_stmt_786_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_554/if_stmt_786_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_554/entry_forx_xend
      -- CP-element group 76: 	 branch_block_stmt_554/entry_forx_xend_PhiReq/$entry
      -- CP-element group 76: 	 branch_block_stmt_554/entry_forx_xend_PhiReq/phi_stmt_1058/$entry
      -- CP-element group 76: 	 branch_block_stmt_554/entry_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_sources/$entry
      -- 
    else_choice_transition_2382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_786_branch_ack_0, ack => convolution3D_CP_1767_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_806_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_806_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_806_Sample/ra
      -- 
    ra_2396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_806_inst_ack_0, ack => convolution3D_CP_1767_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	86 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_806_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_806_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_806_Update/ca
      -- 
    ca_2401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_806_inst_ack_1, ack => convolution3D_CP_1767_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	75 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_822_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_822_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_822_Sample/ra
      -- 
    ra_2410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_822_inst_ack_0, ack => convolution3D_CP_1767_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	75 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_822_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_822_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_822_Update/ca
      -- 
    ca_2415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_822_inst_ack_1, ack => convolution3D_CP_1767_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_831_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_831_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_831_Sample/ra
      -- 
    ra_2424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_831_inst_ack_0, ack => convolution3D_CP_1767_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	75 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_831_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_831_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_831_Update/ca
      -- 
    ca_2429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_831_inst_ack_1, ack => convolution3D_CP_1767_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_841_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_841_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_841_Sample/rr
      -- 
    rr_2437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(83), ack => type_cast_841_inst_req_0); -- 
    convolution3D_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(80) & convolution3D_CP_1767_elements(82);
      gj_convolution3D_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_841_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_841_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_841_Sample/ra
      -- 
    ra_2438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_841_inst_ack_0, ack => convolution3D_CP_1767_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	75 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_841_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_841_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/type_cast_841_Update/ca
      -- 
    ca_2443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_841_inst_ack_1, ack => convolution3D_CP_1767_elements(85)); -- 
    -- CP-element group 86:  join  transition  place  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	78 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	299 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861__exit__
      -- CP-element group 86: 	 branch_block_stmt_554/bbx_xnph369_forx_xbody
      -- CP-element group 86: 	 branch_block_stmt_554/assign_stmt_797_to_assign_stmt_861/$exit
      -- CP-element group 86: 	 branch_block_stmt_554/bbx_xnph369_forx_xbody_PhiReq/$entry
      -- CP-element group 86: 	 branch_block_stmt_554/bbx_xnph369_forx_xbody_PhiReq/phi_stmt_864/$entry
      -- CP-element group 86: 	 branch_block_stmt_554/bbx_xnph369_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_sources/$entry
      -- 
    convolution3D_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(78) & convolution3D_CP_1767_elements(85);
      gj_convolution3D_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	304 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	126 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_final_index_sum_regn_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_final_index_sum_regn_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_final_index_sum_regn_sample_complete
      -- 
    ack_2472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_876_index_offset_ack_0, ack => convolution3D_CP_1767_elements(87)); -- 
    -- CP-element group 88:  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	304 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (11) 
      -- CP-element group 88: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_base_plus_offset/sum_rename_req
      -- CP-element group 88: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_base_plus_offset/$entry
      -- CP-element group 88: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/addr_of_877_request/req
      -- CP-element group 88: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_base_plus_offset/$exit
      -- CP-element group 88: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/addr_of_877_request/$entry
      -- CP-element group 88: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_base_plus_offset/sum_rename_ack
      -- CP-element group 88: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_final_index_sum_regn_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_final_index_sum_regn_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/addr_of_877_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_root_address_calculated
      -- CP-element group 88: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_offset_calculated
      -- 
    ack_2477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_876_index_offset_ack_1, ack => convolution3D_CP_1767_elements(88)); -- 
    req_2486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(88), ack => addr_of_877_final_reg_req_0); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/addr_of_877_request/$exit
      -- CP-element group 89: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/addr_of_877_request/ack
      -- CP-element group 89: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/addr_of_877_sample_completed_
      -- 
    ack_2487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_877_final_reg_ack_0, ack => convolution3D_CP_1767_elements(89)); -- 
    -- CP-element group 90:  fork  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	304 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	123 
    -- CP-element group 90:  members (19) 
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/addr_of_877_complete/$exit
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_word_addrgen/root_register_ack
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_word_addrgen/root_register_req
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_word_addrgen/$exit
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_word_addrgen/$entry
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_base_plus_offset/sum_rename_ack
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_base_plus_offset/sum_rename_req
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_base_plus_offset/$exit
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_base_plus_offset/$entry
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_base_addr_resize/base_resize_ack
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_base_addr_resize/base_resize_req
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_base_addr_resize/$exit
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_base_addr_resize/$entry
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_base_address_resized
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_root_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_word_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_base_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/addr_of_877_complete/ack
      -- CP-element group 90: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/addr_of_877_update_completed_
      -- 
    ack_2492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_877_final_reg_ack_1, ack => convolution3D_CP_1767_elements(90)); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	304 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_880_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_880_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_880_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_880_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_880_update_start_
      -- CP-element group 91: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_880_sample_completed_
      -- 
    ra_2501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_880_inst_ack_0, ack => convolution3D_CP_1767_elements(91)); -- 
    cr_2505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(91), ack => RPIPE_maxpool_input_pipe_880_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92: 	95 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_893_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_893_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_884_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_893_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_884_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_884_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_880_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_880_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_880_update_completed_
      -- 
    ca_2506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_880_inst_ack_1, ack => convolution3D_CP_1767_elements(92)); -- 
    rr_2514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(92), ack => type_cast_884_inst_req_0); -- 
    rr_2528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(92), ack => RPIPE_maxpool_input_pipe_893_inst_req_0); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_884_Sample/ra
      -- CP-element group 93: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_884_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_884_sample_completed_
      -- 
    ra_2515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_884_inst_ack_0, ack => convolution3D_CP_1767_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	304 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	123 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_884_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_884_Update/ca
      -- CP-element group 94: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_884_update_completed_
      -- 
    ca_2520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_884_inst_ack_1, ack => convolution3D_CP_1767_elements(94)); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	92 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_893_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_893_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_893_update_start_
      -- CP-element group 95: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_893_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_893_Update/cr
      -- CP-element group 95: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_893_Update/$entry
      -- 
    ra_2529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_893_inst_ack_0, ack => convolution3D_CP_1767_elements(95)); -- 
    cr_2533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(95), ack => RPIPE_maxpool_input_pipe_893_inst_req_1); -- 
    -- CP-element group 96:  fork  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96: 	99 
    -- CP-element group 96:  members (9) 
      -- CP-element group 96: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_893_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_911_Sample/rr
      -- CP-element group 96: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_911_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_911_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_897_Sample/rr
      -- CP-element group 96: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_897_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_897_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_893_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_893_Update/$exit
      -- 
    ca_2534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_893_inst_ack_1, ack => convolution3D_CP_1767_elements(96)); -- 
    rr_2542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(96), ack => type_cast_897_inst_req_0); -- 
    rr_2556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(96), ack => RPIPE_maxpool_input_pipe_911_inst_req_0); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_897_Sample/ra
      -- CP-element group 97: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_897_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_897_sample_completed_
      -- 
    ra_2543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_897_inst_ack_0, ack => convolution3D_CP_1767_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	304 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	123 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_897_Update/ca
      -- CP-element group 98: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_897_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_897_update_completed_
      -- 
    ca_2548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_897_inst_ack_1, ack => convolution3D_CP_1767_elements(98)); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	96 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_911_Update/cr
      -- CP-element group 99: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_911_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_911_Sample/ra
      -- CP-element group 99: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_911_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_911_update_start_
      -- CP-element group 99: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_911_sample_completed_
      -- 
    ra_2557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_911_inst_ack_0, ack => convolution3D_CP_1767_elements(99)); -- 
    cr_2561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(99), ack => RPIPE_maxpool_input_pipe_911_inst_req_1); -- 
    -- CP-element group 100:  fork  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100: 	103 
    -- CP-element group 100:  members (9) 
      -- CP-element group 100: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_929_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_915_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_929_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_929_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_915_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_915_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_911_Update/ca
      -- CP-element group 100: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_911_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_911_update_completed_
      -- 
    ca_2562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_911_inst_ack_1, ack => convolution3D_CP_1767_elements(100)); -- 
    rr_2570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(100), ack => type_cast_915_inst_req_0); -- 
    rr_2584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(100), ack => RPIPE_maxpool_input_pipe_929_inst_req_0); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_915_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_915_Sample/ra
      -- CP-element group 101: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_915_sample_completed_
      -- 
    ra_2571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_915_inst_ack_0, ack => convolution3D_CP_1767_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	304 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	123 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_915_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_915_Update/ca
      -- CP-element group 102: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_915_update_completed_
      -- 
    ca_2576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_915_inst_ack_1, ack => convolution3D_CP_1767_elements(102)); -- 
    -- CP-element group 103:  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	100 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (6) 
      -- CP-element group 103: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_929_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_929_Update/cr
      -- CP-element group 103: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_929_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_929_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_929_update_start_
      -- CP-element group 103: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_929_Update/$entry
      -- 
    ra_2585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_929_inst_ack_0, ack => convolution3D_CP_1767_elements(103)); -- 
    cr_2589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(103), ack => RPIPE_maxpool_input_pipe_929_inst_req_1); -- 
    -- CP-element group 104:  fork  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	107 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (9) 
      -- CP-element group 104: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_933_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_929_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_933_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_929_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_929_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_933_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_947_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_947_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_947_sample_start_
      -- 
    ca_2590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_929_inst_ack_1, ack => convolution3D_CP_1767_elements(104)); -- 
    rr_2612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(104), ack => RPIPE_maxpool_input_pipe_947_inst_req_0); -- 
    rr_2598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(104), ack => type_cast_933_inst_req_0); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_933_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_933_Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_933_sample_completed_
      -- 
    ra_2599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_933_inst_ack_0, ack => convolution3D_CP_1767_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	304 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	123 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_933_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_933_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_933_Update/ca
      -- 
    ca_2604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_933_inst_ack_1, ack => convolution3D_CP_1767_elements(106)); -- 
    -- CP-element group 107:  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	104 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (6) 
      -- CP-element group 107: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_947_Update/cr
      -- CP-element group 107: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_947_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_947_Sample/ra
      -- CP-element group 107: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_947_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_947_update_start_
      -- CP-element group 107: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_947_sample_completed_
      -- 
    ra_2613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_947_inst_ack_0, ack => convolution3D_CP_1767_elements(107)); -- 
    cr_2617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(107), ack => RPIPE_maxpool_input_pipe_947_inst_req_1); -- 
    -- CP-element group 108:  fork  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108: 	111 
    -- CP-element group 108:  members (9) 
      -- CP-element group 108: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_965_Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_965_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_965_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_951_Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_951_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_951_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_947_Update/ca
      -- CP-element group 108: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_947_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_947_update_completed_
      -- 
    ca_2618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_947_inst_ack_1, ack => convolution3D_CP_1767_elements(108)); -- 
    rr_2626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(108), ack => type_cast_951_inst_req_0); -- 
    rr_2640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(108), ack => RPIPE_maxpool_input_pipe_965_inst_req_0); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_951_Sample/ra
      -- CP-element group 109: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_951_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_951_sample_completed_
      -- 
    ra_2627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_951_inst_ack_0, ack => convolution3D_CP_1767_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	304 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	123 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_951_Update/ca
      -- CP-element group 110: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_951_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_951_update_completed_
      -- 
    ca_2632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_951_inst_ack_1, ack => convolution3D_CP_1767_elements(110)); -- 
    -- CP-element group 111:  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	108 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (6) 
      -- CP-element group 111: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_965_Update/cr
      -- CP-element group 111: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_965_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_965_Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_965_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_965_update_start_
      -- CP-element group 111: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_965_sample_completed_
      -- 
    ra_2641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_965_inst_ack_0, ack => convolution3D_CP_1767_elements(111)); -- 
    cr_2645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(111), ack => RPIPE_maxpool_input_pipe_965_inst_req_1); -- 
    -- CP-element group 112:  fork  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	115 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_983_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_983_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_969_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_969_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_969_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_965_Update/ca
      -- CP-element group 112: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_965_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_965_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_983_Sample/rr
      -- 
    ca_2646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_965_inst_ack_1, ack => convolution3D_CP_1767_elements(112)); -- 
    rr_2654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(112), ack => type_cast_969_inst_req_0); -- 
    rr_2668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(112), ack => RPIPE_maxpool_input_pipe_983_inst_req_0); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_969_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_969_Sample/ra
      -- CP-element group 113: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_969_Sample/$exit
      -- 
    ra_2655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_969_inst_ack_0, ack => convolution3D_CP_1767_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	304 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	123 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_969_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_969_Update/ca
      -- CP-element group 114: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_969_update_completed_
      -- 
    ca_2660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_969_inst_ack_1, ack => convolution3D_CP_1767_elements(114)); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	112 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_983_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_983_update_start_
      -- CP-element group 115: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_983_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_983_Update/cr
      -- CP-element group 115: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_983_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_983_Sample/ra
      -- 
    ra_2669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_983_inst_ack_0, ack => convolution3D_CP_1767_elements(115)); -- 
    cr_2673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(115), ack => RPIPE_maxpool_input_pipe_983_inst_req_1); -- 
    -- CP-element group 116:  fork  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	119 
    -- CP-element group 116:  members (9) 
      -- CP-element group 116: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_1001_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_1001_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_983_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_1001_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_987_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_987_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_987_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_983_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_983_Update/$exit
      -- 
    ca_2674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_983_inst_ack_1, ack => convolution3D_CP_1767_elements(116)); -- 
    rr_2682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(116), ack => type_cast_987_inst_req_0); -- 
    rr_2696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(116), ack => RPIPE_maxpool_input_pipe_1001_inst_req_0); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_987_Sample/ra
      -- CP-element group 117: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_987_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_987_sample_completed_
      -- 
    ra_2683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_987_inst_ack_0, ack => convolution3D_CP_1767_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	304 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	123 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_987_Update/ca
      -- CP-element group 118: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_987_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_987_update_completed_
      -- 
    ca_2688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_987_inst_ack_1, ack => convolution3D_CP_1767_elements(118)); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	116 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (6) 
      -- CP-element group 119: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_1001_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_1001_Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_1001_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_1001_Update/cr
      -- CP-element group 119: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_1001_update_start_
      -- CP-element group 119: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_1001_sample_completed_
      -- 
    ra_2697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1001_inst_ack_0, ack => convolution3D_CP_1767_elements(119)); -- 
    cr_2701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(119), ack => RPIPE_maxpool_input_pipe_1001_inst_req_1); -- 
    -- CP-element group 120:  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (6) 
      -- CP-element group 120: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_1001_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_1005_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_1001_Update/ca
      -- CP-element group 120: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_1001_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_1005_Sample/rr
      -- CP-element group 120: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_1005_Sample/$entry
      -- 
    ca_2702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1001_inst_ack_1, ack => convolution3D_CP_1767_elements(120)); -- 
    rr_2710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(120), ack => type_cast_1005_inst_req_0); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_1005_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_1005_Sample/ra
      -- CP-element group 121: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_1005_Sample/$exit
      -- 
    ra_2711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1005_inst_ack_0, ack => convolution3D_CP_1767_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	304 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_1005_Update/ca
      -- CP-element group 122: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_1005_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_1005_update_completed_
      -- 
    ca_2716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1005_inst_ack_1, ack => convolution3D_CP_1767_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	106 
    -- CP-element group 123: 	110 
    -- CP-element group 123: 	118 
    -- CP-element group 123: 	122 
    -- CP-element group 123: 	114 
    -- CP-element group 123: 	90 
    -- CP-element group 123: 	94 
    -- CP-element group 123: 	98 
    -- CP-element group 123: 	102 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (9) 
      -- CP-element group 123: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Sample/word_access_start/word_0/rr
      -- CP-element group 123: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Sample/ptr_deref_1013_Split/$entry
      -- CP-element group 123: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Sample/word_access_start/word_0/$entry
      -- CP-element group 123: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Sample/ptr_deref_1013_Split/$exit
      -- CP-element group 123: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Sample/word_access_start/$entry
      -- CP-element group 123: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Sample/ptr_deref_1013_Split/split_ack
      -- CP-element group 123: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Sample/ptr_deref_1013_Split/split_req
      -- CP-element group 123: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_sample_start_
      -- 
    rr_2754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(123), ack => ptr_deref_1013_store_0_req_0); -- 
    convolution3D_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(106) & convolution3D_CP_1767_elements(110) & convolution3D_CP_1767_elements(118) & convolution3D_CP_1767_elements(122) & convolution3D_CP_1767_elements(114) & convolution3D_CP_1767_elements(90) & convolution3D_CP_1767_elements(94) & convolution3D_CP_1767_elements(98) & convolution3D_CP_1767_elements(102);
      gj_convolution3D_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Sample/word_access_start/$exit
      -- CP-element group 124: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Sample/word_access_start/word_0/$exit
      -- CP-element group 124: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Sample/word_access_start/word_0/ra
      -- CP-element group 124: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_sample_completed_
      -- 
    ra_2755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1013_store_0_ack_0, ack => convolution3D_CP_1767_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	304 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Update/word_access_complete/word_0/ca
      -- CP-element group 125: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Update/word_access_complete/word_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Update/word_access_complete/$exit
      -- CP-element group 125: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_update_completed_
      -- 
    ca_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1013_store_0_ack_1, ack => convolution3D_CP_1767_elements(125)); -- 
    -- CP-element group 126:  branch  join  transition  place  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: 	87 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (10) 
      -- CP-element group 126: 	 branch_block_stmt_554/if_stmt_1027_dead_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026__exit__
      -- CP-element group 126: 	 branch_block_stmt_554/if_stmt_1027__entry__
      -- CP-element group 126: 	 branch_block_stmt_554/if_stmt_1027_eval_test/$entry
      -- CP-element group 126: 	 branch_block_stmt_554/if_stmt_1027_eval_test/branch_req
      -- CP-element group 126: 	 branch_block_stmt_554/if_stmt_1027_eval_test/$exit
      -- CP-element group 126: 	 branch_block_stmt_554/R_exitcond28_1028_place
      -- CP-element group 126: 	 branch_block_stmt_554/if_stmt_1027_else_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_554/if_stmt_1027_if_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/$exit
      -- 
    branch_req_2774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(126), ack => if_stmt_1027_branch_req_0); -- 
    convolution3D_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(125) & convolution3D_CP_1767_elements(87);
      gj_convolution3D_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	306 
    -- CP-element group 127: 	307 
    -- CP-element group 127:  members (24) 
      -- CP-element group 127: 	 branch_block_stmt_554/merge_stmt_1033__exit__
      -- CP-element group 127: 	 branch_block_stmt_554/assign_stmt_1040_to_assign_stmt_1055__entry__
      -- CP-element group 127: 	 branch_block_stmt_554/assign_stmt_1040_to_assign_stmt_1055__exit__
      -- CP-element group 127: 	 branch_block_stmt_554/forx_xbody_forx_xcondx_xforx_xend_crit_edge
      -- CP-element group 127: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend
      -- CP-element group 127: 	 branch_block_stmt_554/assign_stmt_1040_to_assign_stmt_1055/$exit
      -- CP-element group 127: 	 branch_block_stmt_554/assign_stmt_1040_to_assign_stmt_1055/$entry
      -- CP-element group 127: 	 branch_block_stmt_554/if_stmt_1027_if_link/if_choice_transition
      -- CP-element group 127: 	 branch_block_stmt_554/if_stmt_1027_if_link/$exit
      -- CP-element group 127: 	 branch_block_stmt_554/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_554/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$exit
      -- CP-element group 127: 	 branch_block_stmt_554/merge_stmt_1033_PhiReqMerge
      -- CP-element group 127: 	 branch_block_stmt_554/merge_stmt_1033_PhiAck/$entry
      -- CP-element group 127: 	 branch_block_stmt_554/merge_stmt_1033_PhiAck/$exit
      -- CP-element group 127: 	 branch_block_stmt_554/merge_stmt_1033_PhiAck/dummy
      -- CP-element group 127: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1058/$entry
      -- CP-element group 127: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_sources/$entry
      -- CP-element group 127: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_sources/type_cast_1061/$entry
      -- CP-element group 127: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_sources/type_cast_1061/SplitProtocol/$entry
      -- CP-element group 127: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_sources/type_cast_1061/SplitProtocol/Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_sources/type_cast_1061/SplitProtocol/Sample/rr
      -- CP-element group 127: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_sources/type_cast_1061/SplitProtocol/Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_sources/type_cast_1061/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1027_branch_ack_1, ack => convolution3D_CP_1767_elements(127)); -- 
    rr_4196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(127), ack => type_cast_1061_inst_req_0); -- 
    cr_4201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(127), ack => type_cast_1061_inst_req_1); -- 
    -- CP-element group 128:  fork  transition  place  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	300 
    -- CP-element group 128: 	301 
    -- CP-element group 128:  members (12) 
      -- CP-element group 128: 	 branch_block_stmt_554/forx_xbody_forx_xbody
      -- CP-element group 128: 	 branch_block_stmt_554/if_stmt_1027_else_link/else_choice_transition
      -- CP-element group 128: 	 branch_block_stmt_554/if_stmt_1027_else_link/$exit
      -- CP-element group 128: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 128: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/phi_stmt_864/$entry
      -- CP-element group 128: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_sources/$entry
      -- CP-element group 128: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_sources/type_cast_870/$entry
      -- CP-element group 128: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_sources/type_cast_870/SplitProtocol/$entry
      -- CP-element group 128: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_sources/type_cast_870/SplitProtocol/Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_sources/type_cast_870/SplitProtocol/Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_sources/type_cast_870/SplitProtocol/Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_sources/type_cast_870/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1027_branch_ack_0, ack => convolution3D_CP_1767_elements(128)); -- 
    rr_4142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(128), ack => type_cast_870_inst_req_0); -- 
    cr_4147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(128), ack => type_cast_870_inst_req_1); -- 
    -- CP-element group 129:  transition  place  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	310 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	329 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_554/if_stmt_1078_if_link/$exit
      -- CP-element group 129: 	 branch_block_stmt_554/forx_xend_ifx_xend
      -- CP-element group 129: 	 branch_block_stmt_554/if_stmt_1078_if_link/if_choice_transition
      -- CP-element group 129: 	 branch_block_stmt_554/forx_xend_ifx_xend_PhiReq/$entry
      -- CP-element group 129: 	 branch_block_stmt_554/forx_xend_ifx_xend_PhiReq/$exit
      -- 
    if_choice_transition_2804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1078_branch_ack_1, ack => convolution3D_CP_1767_elements(129)); -- 
    -- CP-element group 130:  merge  fork  transition  place  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	310 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	311 
    -- CP-element group 130: 	312 
    -- CP-element group 130:  members (20) 
      -- CP-element group 130: 	 branch_block_stmt_554/assign_stmt_1090_to_assign_stmt_1096/$entry
      -- CP-element group 130: 	 branch_block_stmt_554/if_stmt_1078_else_link/else_choice_transition
      -- CP-element group 130: 	 branch_block_stmt_554/bbx_xnphx_xi_forx_xbodyx_xi
      -- CP-element group 130: 	 branch_block_stmt_554/assign_stmt_1090_to_assign_stmt_1096__exit__
      -- CP-element group 130: 	 branch_block_stmt_554/assign_stmt_1090_to_assign_stmt_1096__entry__
      -- CP-element group 130: 	 branch_block_stmt_554/merge_stmt_1084__exit__
      -- CP-element group 130: 	 branch_block_stmt_554/if_stmt_1078_else_link/$exit
      -- CP-element group 130: 	 branch_block_stmt_554/forx_xend_bbx_xnphx_xi
      -- CP-element group 130: 	 branch_block_stmt_554/assign_stmt_1090_to_assign_stmt_1096/$exit
      -- CP-element group 130: 	 branch_block_stmt_554/forx_xend_bbx_xnphx_xi_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_554/forx_xend_bbx_xnphx_xi_PhiReq/$exit
      -- CP-element group 130: 	 branch_block_stmt_554/merge_stmt_1084_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_554/merge_stmt_1084_PhiAck/$entry
      -- CP-element group 130: 	 branch_block_stmt_554/merge_stmt_1084_PhiAck/$exit
      -- CP-element group 130: 	 branch_block_stmt_554/merge_stmt_1084_PhiAck/dummy
      -- CP-element group 130: 	 branch_block_stmt_554/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_554/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/$entry
      -- CP-element group 130: 	 branch_block_stmt_554/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_554/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/$entry
      -- CP-element group 130: 	 branch_block_stmt_554/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/$entry
      -- 
    else_choice_transition_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1078_branch_ack_0, ack => convolution3D_CP_1767_elements(130)); -- 
    -- CP-element group 131:  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	324 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (6) 
      -- CP-element group 131: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/RPIPE_maxpool_input_pipe_1127_Update/cr
      -- CP-element group 131: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/RPIPE_maxpool_input_pipe_1127_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/RPIPE_maxpool_input_pipe_1127_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/RPIPE_maxpool_input_pipe_1127_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/RPIPE_maxpool_input_pipe_1127_update_start_
      -- CP-element group 131: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/RPIPE_maxpool_input_pipe_1127_sample_completed_
      -- 
    ra_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1127_inst_ack_0, ack => convolution3D_CP_1767_elements(131)); -- 
    cr_2829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(131), ack => RPIPE_maxpool_input_pipe_1127_inst_req_1); -- 
    -- CP-element group 132:  transition  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (6) 
      -- CP-element group 132: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1131_Sample/rr
      -- CP-element group 132: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1131_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1131_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/RPIPE_maxpool_input_pipe_1127_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/RPIPE_maxpool_input_pipe_1127_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/RPIPE_maxpool_input_pipe_1127_update_completed_
      -- 
    ca_2830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1127_inst_ack_1, ack => convolution3D_CP_1767_elements(132)); -- 
    rr_2838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(132), ack => type_cast_1131_inst_req_0); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1131_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1131_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1131_sample_completed_
      -- 
    ra_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1131_inst_ack_0, ack => convolution3D_CP_1767_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	324 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1131_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1131_Update/ca
      -- CP-element group 134: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1131_update_completed_
      -- 
    ca_2844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1131_inst_ack_1, ack => convolution3D_CP_1767_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	324 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1146_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1146_Sample/ra
      -- CP-element group 135: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1146_Sample/$exit
      -- 
    ra_2853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1146_inst_ack_0, ack => convolution3D_CP_1767_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	324 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1146_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1146_Update/ca
      -- CP-element group 136: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1146_Update/$exit
      -- 
    ca_2858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1146_inst_ack_1, ack => convolution3D_CP_1767_elements(136)); -- 
    -- CP-element group 137:  branch  join  transition  place  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (10) 
      -- CP-element group 137: 	 branch_block_stmt_554/if_stmt_1153_eval_test/$exit
      -- CP-element group 137: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152__exit__
      -- CP-element group 137: 	 branch_block_stmt_554/if_stmt_1153__entry__
      -- CP-element group 137: 	 branch_block_stmt_554/R_cmpx_xi_1154_place
      -- CP-element group 137: 	 branch_block_stmt_554/if_stmt_1153_eval_test/$entry
      -- CP-element group 137: 	 branch_block_stmt_554/if_stmt_1153_eval_test/branch_req
      -- CP-element group 137: 	 branch_block_stmt_554/if_stmt_1153_if_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_554/if_stmt_1153_dead_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_554/if_stmt_1153_else_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/$exit
      -- 
    branch_req_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(137), ack => if_stmt_1153_branch_req_0); -- 
    convolution3D_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(134) & convolution3D_CP_1767_elements(136);
      gj_convolution3D_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  place  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	314 
    -- CP-element group 138: 	315 
    -- CP-element group 138: 	317 
    -- CP-element group 138: 	318 
    -- CP-element group 138:  members (20) 
      -- CP-element group 138: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi
      -- CP-element group 138: 	 branch_block_stmt_554/if_stmt_1153_if_link/if_choice_transition
      -- CP-element group 138: 	 branch_block_stmt_554/if_stmt_1153_if_link/$exit
      -- CP-element group 138: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 138: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/$entry
      -- CP-element group 138: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_sources/$entry
      -- CP-element group 138: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_sources/type_cast_1105/$entry
      -- CP-element group 138: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_sources/type_cast_1105/SplitProtocol/$entry
      -- CP-element group 138: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_sources/type_cast_1105/SplitProtocol/Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_sources/type_cast_1105/SplitProtocol/Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_sources/type_cast_1105/SplitProtocol/Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_sources/type_cast_1105/SplitProtocol/Update/cr
      -- CP-element group 138: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/$entry
      -- CP-element group 138: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/$entry
      -- CP-element group 138: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/$entry
      -- CP-element group 138: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/$entry
      -- CP-element group 138: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1153_branch_ack_1, ack => convolution3D_CP_1767_elements(138)); -- 
    rr_4258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(138), ack => type_cast_1105_inst_req_0); -- 
    cr_4263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(138), ack => type_cast_1105_inst_req_1); -- 
    rr_4281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(138), ack => type_cast_1112_inst_req_0); -- 
    cr_4286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(138), ack => type_cast_1112_inst_req_1); -- 
    -- CP-element group 139:  fork  transition  place  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	325 
    -- CP-element group 139: 	326 
    -- CP-element group 139:  members (12) 
      -- CP-element group 139: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit
      -- CP-element group 139: 	 branch_block_stmt_554/if_stmt_1153_else_link/else_choice_transition
      -- CP-element group 139: 	 branch_block_stmt_554/if_stmt_1153_else_link/$exit
      -- CP-element group 139: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 139: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1160/$entry
      -- CP-element group 139: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1160/phi_stmt_1160_sources/$entry
      -- CP-element group 139: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1160/phi_stmt_1160_sources/type_cast_1163/$entry
      -- CP-element group 139: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1160/phi_stmt_1160_sources/type_cast_1163/SplitProtocol/$entry
      -- CP-element group 139: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1160/phi_stmt_1160_sources/type_cast_1163/SplitProtocol/Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1160/phi_stmt_1160_sources/type_cast_1163/SplitProtocol/Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1160/phi_stmt_1160_sources/type_cast_1163/SplitProtocol/Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1160/phi_stmt_1160_sources/type_cast_1163/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1153_branch_ack_0, ack => convolution3D_CP_1767_elements(139)); -- 
    rr_4317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(139), ack => type_cast_1163_inst_req_0); -- 
    cr_4322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(139), ack => type_cast_1163_inst_req_1); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	328 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	146 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_final_index_sum_regn_sample_complete
      -- CP-element group 140: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_final_index_sum_regn_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_final_index_sum_regn_Sample/ack
      -- 
    ack_2906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1192_index_offset_ack_0, ack => convolution3D_CP_1767_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	328 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (11) 
      -- CP-element group 141: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_root_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/addr_of_1193_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_offset_calculated
      -- CP-element group 141: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_final_index_sum_regn_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_final_index_sum_regn_Update/ack
      -- CP-element group 141: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_base_plus_offset/$entry
      -- CP-element group 141: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_base_plus_offset/$exit
      -- CP-element group 141: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_base_plus_offset/sum_rename_req
      -- CP-element group 141: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_base_plus_offset/sum_rename_ack
      -- CP-element group 141: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/addr_of_1193_request/$entry
      -- CP-element group 141: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/addr_of_1193_request/req
      -- 
    ack_2911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1192_index_offset_ack_1, ack => convolution3D_CP_1767_elements(141)); -- 
    req_2920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(141), ack => addr_of_1193_final_reg_req_0); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/addr_of_1193_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/addr_of_1193_request/$exit
      -- CP-element group 142: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/addr_of_1193_request/ack
      -- 
    ack_2921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1193_final_reg_ack_0, ack => convolution3D_CP_1767_elements(142)); -- 
    -- CP-element group 143:  join  fork  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	328 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (28) 
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/addr_of_1193_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/addr_of_1193_complete/$exit
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/addr_of_1193_complete/ack
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_base_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_word_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_root_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_base_address_resized
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_base_addr_resize/$entry
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_base_addr_resize/$exit
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_base_addr_resize/base_resize_req
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_base_addr_resize/base_resize_ack
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_base_plus_offset/$entry
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_base_plus_offset/$exit
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_base_plus_offset/sum_rename_req
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_base_plus_offset/sum_rename_ack
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_word_addrgen/$entry
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_word_addrgen/$exit
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_word_addrgen/root_register_req
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_word_addrgen/root_register_ack
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Sample/ptr_deref_1196_Split/$entry
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Sample/ptr_deref_1196_Split/$exit
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Sample/ptr_deref_1196_Split/split_req
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Sample/ptr_deref_1196_Split/split_ack
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Sample/word_access_start/$entry
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Sample/word_access_start/word_0/$entry
      -- CP-element group 143: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Sample/word_access_start/word_0/rr
      -- 
    ack_2926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1193_final_reg_ack_1, ack => convolution3D_CP_1767_elements(143)); -- 
    rr_2964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(143), ack => ptr_deref_1196_store_0_req_0); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Sample/word_access_start/$exit
      -- CP-element group 144: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Sample/word_access_start/word_0/$exit
      -- CP-element group 144: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Sample/word_access_start/word_0/ra
      -- 
    ra_2965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1196_store_0_ack_0, ack => convolution3D_CP_1767_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	328 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (5) 
      -- CP-element group 145: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Update/word_access_complete/$exit
      -- CP-element group 145: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Update/word_access_complete/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Update/word_access_complete/word_0/ca
      -- 
    ca_2976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1196_store_0_ack_1, ack => convolution3D_CP_1767_elements(145)); -- 
    -- CP-element group 146:  join  transition  place  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: 	140 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	329 
    -- CP-element group 146:  members (5) 
      -- CP-element group 146: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198__exit__
      -- CP-element group 146: 	 branch_block_stmt_554/getRemainingElementsx_xexit_ifx_xend
      -- CP-element group 146: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/$exit
      -- CP-element group 146: 	 branch_block_stmt_554/getRemainingElementsx_xexit_ifx_xend_PhiReq/$entry
      -- CP-element group 146: 	 branch_block_stmt_554/getRemainingElementsx_xexit_ifx_xend_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(145) & convolution3D_CP_1767_elements(140);
      gj_convolution3D_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	329 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1203_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1203_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1203_Sample/ra
      -- 
    ra_2988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1203_inst_ack_0, ack => convolution3D_CP_1767_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	329 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	153 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1203_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1203_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1203_Update/ca
      -- 
    ca_2993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1203_inst_ack_1, ack => convolution3D_CP_1767_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	329 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1207_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1207_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1207_Sample/ra
      -- 
    ra_3002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1207_inst_ack_0, ack => convolution3D_CP_1767_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	329 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	153 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1207_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1207_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1207_Update/ca
      -- 
    ca_3007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1207_inst_ack_1, ack => convolution3D_CP_1767_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	329 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1211_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1211_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1211_Sample/ra
      -- 
    ra_3016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1211_inst_ack_0, ack => convolution3D_CP_1767_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	329 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1211_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1211_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1211_Update/ca
      -- 
    ca_3021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1211_inst_ack_1, ack => convolution3D_CP_1767_elements(152)); -- 
    -- CP-element group 153:  branch  join  transition  place  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: 	150 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (10) 
      -- CP-element group 153: 	 branch_block_stmt_554/if_stmt_1249__entry__
      -- CP-element group 153: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248__exit__
      -- CP-element group 153: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/$exit
      -- CP-element group 153: 	 branch_block_stmt_554/if_stmt_1249_dead_link/$entry
      -- CP-element group 153: 	 branch_block_stmt_554/if_stmt_1249_eval_test/$entry
      -- CP-element group 153: 	 branch_block_stmt_554/if_stmt_1249_eval_test/$exit
      -- CP-element group 153: 	 branch_block_stmt_554/if_stmt_1249_eval_test/branch_req
      -- CP-element group 153: 	 branch_block_stmt_554/R_cmp161363_1250_place
      -- CP-element group 153: 	 branch_block_stmt_554/if_stmt_1249_if_link/$entry
      -- CP-element group 153: 	 branch_block_stmt_554/if_stmt_1249_else_link/$entry
      -- 
    branch_req_3029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(153), ack => if_stmt_1249_branch_req_0); -- 
    convolution3D_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(148) & convolution3D_CP_1767_elements(150) & convolution3D_CP_1767_elements(152);
      gj_convolution3D_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	160 
    -- CP-element group 154: 	161 
    -- CP-element group 154: 	164 
    -- CP-element group 154: 	158 
    -- CP-element group 154: 	159 
    -- CP-element group 154: 	156 
    -- CP-element group 154: 	157 
    -- CP-element group 154: 	166 
    -- CP-element group 154:  members (36) 
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322__entry__
      -- CP-element group 154: 	 branch_block_stmt_554/merge_stmt_1255__exit__
      -- CP-element group 154: 	 branch_block_stmt_554/if_stmt_1249_if_link/$exit
      -- CP-element group 154: 	 branch_block_stmt_554/if_stmt_1249_if_link/if_choice_transition
      -- CP-element group 154: 	 branch_block_stmt_554/ifx_xend_bbx_xnph
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/$entry
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1270_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1270_update_start_
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1270_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1270_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1270_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1270_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1279_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1279_update_start_
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1279_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1279_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1279_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1279_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1288_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1288_update_start_
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1288_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1288_Sample/rr
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1288_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1288_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1297_update_start_
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1297_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1297_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1302_update_start_
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1302_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1302_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_554/ifx_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 154: 	 branch_block_stmt_554/ifx_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 154: 	 branch_block_stmt_554/merge_stmt_1255_PhiReqMerge
      -- CP-element group 154: 	 branch_block_stmt_554/merge_stmt_1255_PhiAck/$entry
      -- CP-element group 154: 	 branch_block_stmt_554/merge_stmt_1255_PhiAck/$exit
      -- CP-element group 154: 	 branch_block_stmt_554/merge_stmt_1255_PhiAck/dummy
      -- 
    if_choice_transition_3034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1249_branch_ack_1, ack => convolution3D_CP_1767_elements(154)); -- 
    rr_3051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(154), ack => type_cast_1270_inst_req_0); -- 
    cr_3056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(154), ack => type_cast_1270_inst_req_1); -- 
    rr_3065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(154), ack => type_cast_1279_inst_req_0); -- 
    cr_3070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(154), ack => type_cast_1279_inst_req_1); -- 
    rr_3079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(154), ack => type_cast_1288_inst_req_0); -- 
    cr_3084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(154), ack => type_cast_1288_inst_req_1); -- 
    cr_3098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(154), ack => type_cast_1297_inst_req_1); -- 
    cr_3112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(154), ack => type_cast_1302_inst_req_1); -- 
    -- CP-element group 155:  transition  place  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	339 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_554/if_stmt_1249_else_link/$exit
      -- CP-element group 155: 	 branch_block_stmt_554/if_stmt_1249_else_link/else_choice_transition
      -- CP-element group 155: 	 branch_block_stmt_554/ifx_xend_forx_xend215
      -- CP-element group 155: 	 branch_block_stmt_554/ifx_xend_forx_xend215_PhiReq/$entry
      -- CP-element group 155: 	 branch_block_stmt_554/ifx_xend_forx_xend215_PhiReq/phi_stmt_1519/$entry
      -- CP-element group 155: 	 branch_block_stmt_554/ifx_xend_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/$entry
      -- 
    else_choice_transition_3038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1249_branch_ack_0, ack => convolution3D_CP_1767_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1270_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1270_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1270_Sample/ra
      -- 
    ra_3052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1270_inst_ack_0, ack => convolution3D_CP_1767_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	154 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	162 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1270_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1270_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1270_Update/ca
      -- 
    ca_3057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1270_inst_ack_1, ack => convolution3D_CP_1767_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	154 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1279_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1279_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1279_Sample/ra
      -- 
    ra_3066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1279_inst_ack_0, ack => convolution3D_CP_1767_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	154 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	162 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1279_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1279_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1279_Update/ca
      -- 
    ca_3071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1279_inst_ack_1, ack => convolution3D_CP_1767_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	154 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1288_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1288_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1288_Sample/ra
      -- 
    ra_3080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1288_inst_ack_0, ack => convolution3D_CP_1767_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	154 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1288_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1288_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1288_Update/ca
      -- 
    ca_3085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1288_inst_ack_1, ack => convolution3D_CP_1767_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: 	159 
    -- CP-element group 162: 	157 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1297_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1297_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1297_Sample/rr
      -- 
    rr_3093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(162), ack => type_cast_1297_inst_req_0); -- 
    convolution3D_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(161) & convolution3D_CP_1767_elements(159) & convolution3D_CP_1767_elements(157);
      gj_convolution3D_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1297_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1297_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1297_Sample/ra
      -- 
    ra_3094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1297_inst_ack_0, ack => convolution3D_CP_1767_elements(163)); -- 
    -- CP-element group 164:  transition  input  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	154 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (6) 
      -- CP-element group 164: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1297_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1297_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1297_Update/ca
      -- CP-element group 164: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1302_sample_start_
      -- CP-element group 164: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1302_Sample/$entry
      -- CP-element group 164: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1302_Sample/rr
      -- 
    ca_3099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1297_inst_ack_1, ack => convolution3D_CP_1767_elements(164)); -- 
    rr_3107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(164), ack => type_cast_1302_inst_req_0); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1302_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1302_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1302_Sample/ra
      -- 
    ra_3108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1302_inst_ack_0, ack => convolution3D_CP_1767_elements(165)); -- 
    -- CP-element group 166:  transition  place  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	154 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	330 
    -- CP-element group 166:  members (9) 
      -- CP-element group 166: 	 branch_block_stmt_554/bbx_xnph_forx_xbody163
      -- CP-element group 166: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322__exit__
      -- CP-element group 166: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/$exit
      -- CP-element group 166: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1302_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1302_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_554/assign_stmt_1261_to_assign_stmt_1322/type_cast_1302_Update/ca
      -- CP-element group 166: 	 branch_block_stmt_554/bbx_xnph_forx_xbody163_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_554/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1325/$entry
      -- CP-element group 166: 	 branch_block_stmt_554/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_sources/$entry
      -- 
    ca_3113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1302_inst_ack_1, ack => convolution3D_CP_1767_elements(166)); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	335 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	206 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_final_index_sum_regn_sample_complete
      -- CP-element group 167: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_final_index_sum_regn_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_final_index_sum_regn_Sample/ack
      -- 
    ack_3142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1337_index_offset_ack_0, ack => convolution3D_CP_1767_elements(167)); -- 
    -- CP-element group 168:  transition  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	335 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (11) 
      -- CP-element group 168: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/addr_of_1338_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_root_address_calculated
      -- CP-element group 168: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_offset_calculated
      -- CP-element group 168: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_final_index_sum_regn_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_final_index_sum_regn_Update/ack
      -- CP-element group 168: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_base_plus_offset/$entry
      -- CP-element group 168: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_base_plus_offset/$exit
      -- CP-element group 168: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_base_plus_offset/sum_rename_req
      -- CP-element group 168: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_base_plus_offset/sum_rename_ack
      -- CP-element group 168: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/addr_of_1338_request/$entry
      -- CP-element group 168: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/addr_of_1338_request/req
      -- 
    ack_3147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1337_index_offset_ack_1, ack => convolution3D_CP_1767_elements(168)); -- 
    req_3156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(168), ack => addr_of_1338_final_reg_req_0); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/addr_of_1338_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/addr_of_1338_request/$exit
      -- CP-element group 169: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/addr_of_1338_request/ack
      -- 
    ack_3157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1338_final_reg_ack_0, ack => convolution3D_CP_1767_elements(169)); -- 
    -- CP-element group 170:  fork  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	335 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	203 
    -- CP-element group 170:  members (19) 
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/addr_of_1338_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/addr_of_1338_complete/$exit
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/addr_of_1338_complete/ack
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_base_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_word_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_root_address_calculated
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_base_address_resized
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_base_addr_resize/$entry
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_base_addr_resize/$exit
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_base_addr_resize/base_resize_req
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_base_addr_resize/base_resize_ack
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_base_plus_offset/$entry
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_base_plus_offset/$exit
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_base_plus_offset/sum_rename_req
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_base_plus_offset/sum_rename_ack
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_word_addrgen/$entry
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_word_addrgen/$exit
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_word_addrgen/root_register_req
      -- CP-element group 170: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_word_addrgen/root_register_ack
      -- 
    ack_3162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1338_final_reg_ack_1, ack => convolution3D_CP_1767_elements(170)); -- 
    -- CP-element group 171:  transition  input  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	335 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (6) 
      -- CP-element group 171: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1341_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1341_update_start_
      -- CP-element group 171: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1341_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1341_Sample/ra
      -- CP-element group 171: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1341_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1341_Update/cr
      -- 
    ra_3171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1341_inst_ack_0, ack => convolution3D_CP_1767_elements(171)); -- 
    cr_3175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(171), ack => RPIPE_maxpool_input_pipe_1341_inst_req_1); -- 
    -- CP-element group 172:  fork  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172: 	175 
    -- CP-element group 172:  members (9) 
      -- CP-element group 172: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1341_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1341_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1341_Update/ca
      -- CP-element group 172: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1345_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1345_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1345_Sample/rr
      -- CP-element group 172: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1354_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1354_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1354_Sample/rr
      -- 
    ca_3176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1341_inst_ack_1, ack => convolution3D_CP_1767_elements(172)); -- 
    rr_3184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(172), ack => type_cast_1345_inst_req_0); -- 
    rr_3198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(172), ack => RPIPE_maxpool_input_pipe_1354_inst_req_0); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1345_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1345_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1345_Sample/ra
      -- 
    ra_3185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1345_inst_ack_0, ack => convolution3D_CP_1767_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	335 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	203 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1345_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1345_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1345_Update/ca
      -- 
    ca_3190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1345_inst_ack_1, ack => convolution3D_CP_1767_elements(174)); -- 
    -- CP-element group 175:  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	172 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (6) 
      -- CP-element group 175: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1354_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1354_update_start_
      -- CP-element group 175: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1354_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1354_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1354_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1354_Update/cr
      -- 
    ra_3199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1354_inst_ack_0, ack => convolution3D_CP_1767_elements(175)); -- 
    cr_3203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(175), ack => RPIPE_maxpool_input_pipe_1354_inst_req_1); -- 
    -- CP-element group 176:  fork  transition  input  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176: 	179 
    -- CP-element group 176:  members (9) 
      -- CP-element group 176: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1354_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1354_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1354_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1358_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1358_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1358_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1372_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1372_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1372_Sample/rr
      -- 
    ca_3204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1354_inst_ack_1, ack => convolution3D_CP_1767_elements(176)); -- 
    rr_3212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(176), ack => type_cast_1358_inst_req_0); -- 
    rr_3226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(176), ack => RPIPE_maxpool_input_pipe_1372_inst_req_0); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1358_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1358_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1358_Sample/ra
      -- 
    ra_3213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1358_inst_ack_0, ack => convolution3D_CP_1767_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	335 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	203 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1358_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1358_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1358_Update/ca
      -- 
    ca_3218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1358_inst_ack_1, ack => convolution3D_CP_1767_elements(178)); -- 
    -- CP-element group 179:  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	176 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1372_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1372_update_start_
      -- CP-element group 179: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1372_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1372_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1372_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1372_Update/cr
      -- 
    ra_3227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1372_inst_ack_0, ack => convolution3D_CP_1767_elements(179)); -- 
    cr_3231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(179), ack => RPIPE_maxpool_input_pipe_1372_inst_req_1); -- 
    -- CP-element group 180:  fork  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: 	183 
    -- CP-element group 180:  members (9) 
      -- CP-element group 180: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1372_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1372_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1372_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1376_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1376_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1376_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1390_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1390_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1390_Sample/rr
      -- 
    ca_3232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1372_inst_ack_1, ack => convolution3D_CP_1767_elements(180)); -- 
    rr_3240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(180), ack => type_cast_1376_inst_req_0); -- 
    rr_3254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(180), ack => RPIPE_maxpool_input_pipe_1390_inst_req_0); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1376_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1376_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1376_Sample/ra
      -- 
    ra_3241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1376_inst_ack_0, ack => convolution3D_CP_1767_elements(181)); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	335 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	203 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1376_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1376_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1376_Update/ca
      -- 
    ca_3246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1376_inst_ack_1, ack => convolution3D_CP_1767_elements(182)); -- 
    -- CP-element group 183:  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	180 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (6) 
      -- CP-element group 183: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1390_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1390_update_start_
      -- CP-element group 183: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1390_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1390_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1390_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1390_Update/cr
      -- 
    ra_3255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1390_inst_ack_0, ack => convolution3D_CP_1767_elements(183)); -- 
    cr_3259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(183), ack => RPIPE_maxpool_input_pipe_1390_inst_req_1); -- 
    -- CP-element group 184:  fork  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	187 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (9) 
      -- CP-element group 184: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1390_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1390_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1390_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1394_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1394_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1394_Sample/rr
      -- CP-element group 184: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1408_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1408_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1408_Sample/rr
      -- 
    ca_3260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1390_inst_ack_1, ack => convolution3D_CP_1767_elements(184)); -- 
    rr_3282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(184), ack => RPIPE_maxpool_input_pipe_1408_inst_req_0); -- 
    rr_3268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(184), ack => type_cast_1394_inst_req_0); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1394_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1394_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1394_Sample/ra
      -- 
    ra_3269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1394_inst_ack_0, ack => convolution3D_CP_1767_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	335 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	203 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1394_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1394_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1394_Update/ca
      -- 
    ca_3274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1394_inst_ack_1, ack => convolution3D_CP_1767_elements(186)); -- 
    -- CP-element group 187:  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	184 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1408_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1408_update_start_
      -- CP-element group 187: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1408_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1408_Sample/ra
      -- CP-element group 187: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1408_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1408_Update/cr
      -- 
    ra_3283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1408_inst_ack_0, ack => convolution3D_CP_1767_elements(187)); -- 
    cr_3287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(187), ack => RPIPE_maxpool_input_pipe_1408_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188: 	191 
    -- CP-element group 188:  members (9) 
      -- CP-element group 188: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1408_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1408_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1408_Update/ca
      -- CP-element group 188: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1412_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1412_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1412_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1426_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1426_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1426_Sample/rr
      -- 
    ca_3288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1408_inst_ack_1, ack => convolution3D_CP_1767_elements(188)); -- 
    rr_3296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(188), ack => type_cast_1412_inst_req_0); -- 
    rr_3310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(188), ack => RPIPE_maxpool_input_pipe_1426_inst_req_0); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1412_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1412_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1412_Sample/ra
      -- 
    ra_3297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1412_inst_ack_0, ack => convolution3D_CP_1767_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	335 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	203 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1412_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1412_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1412_Update/ca
      -- 
    ca_3302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1412_inst_ack_1, ack => convolution3D_CP_1767_elements(190)); -- 
    -- CP-element group 191:  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	188 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (6) 
      -- CP-element group 191: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1426_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1426_update_start_
      -- CP-element group 191: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1426_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1426_Sample/ra
      -- CP-element group 191: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1426_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1426_Update/cr
      -- 
    ra_3311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1426_inst_ack_0, ack => convolution3D_CP_1767_elements(191)); -- 
    cr_3315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(191), ack => RPIPE_maxpool_input_pipe_1426_inst_req_1); -- 
    -- CP-element group 192:  fork  transition  input  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192: 	195 
    -- CP-element group 192:  members (9) 
      -- CP-element group 192: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1426_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1426_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1426_Update/ca
      -- CP-element group 192: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1430_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1430_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1430_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1444_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1444_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1444_Sample/rr
      -- 
    ca_3316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1426_inst_ack_1, ack => convolution3D_CP_1767_elements(192)); -- 
    rr_3324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(192), ack => type_cast_1430_inst_req_0); -- 
    rr_3338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(192), ack => RPIPE_maxpool_input_pipe_1444_inst_req_0); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1430_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1430_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1430_Sample/ra
      -- 
    ra_3325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1430_inst_ack_0, ack => convolution3D_CP_1767_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	335 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	203 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1430_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1430_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1430_Update/ca
      -- 
    ca_3330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1430_inst_ack_1, ack => convolution3D_CP_1767_elements(194)); -- 
    -- CP-element group 195:  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	192 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (6) 
      -- CP-element group 195: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1444_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1444_update_start_
      -- CP-element group 195: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1444_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1444_Sample/ra
      -- CP-element group 195: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1444_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1444_Update/cr
      -- 
    ra_3339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1444_inst_ack_0, ack => convolution3D_CP_1767_elements(195)); -- 
    cr_3343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(195), ack => RPIPE_maxpool_input_pipe_1444_inst_req_1); -- 
    -- CP-element group 196:  fork  transition  input  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196: 	199 
    -- CP-element group 196:  members (9) 
      -- CP-element group 196: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1444_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1444_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1444_Update/ca
      -- CP-element group 196: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1448_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1448_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1448_Sample/rr
      -- CP-element group 196: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1462_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1462_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1462_Sample/rr
      -- 
    ca_3344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1444_inst_ack_1, ack => convolution3D_CP_1767_elements(196)); -- 
    rr_3352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(196), ack => type_cast_1448_inst_req_0); -- 
    rr_3366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(196), ack => RPIPE_maxpool_input_pipe_1462_inst_req_0); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1448_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1448_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1448_Sample/ra
      -- 
    ra_3353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1448_inst_ack_0, ack => convolution3D_CP_1767_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	335 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	203 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1448_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1448_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1448_Update/ca
      -- 
    ca_3358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1448_inst_ack_1, ack => convolution3D_CP_1767_elements(198)); -- 
    -- CP-element group 199:  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	196 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (6) 
      -- CP-element group 199: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1462_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1462_update_start_
      -- CP-element group 199: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1462_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1462_Sample/ra
      -- CP-element group 199: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1462_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1462_Update/cr
      -- 
    ra_3367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1462_inst_ack_0, ack => convolution3D_CP_1767_elements(199)); -- 
    cr_3371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(199), ack => RPIPE_maxpool_input_pipe_1462_inst_req_1); -- 
    -- CP-element group 200:  transition  input  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (6) 
      -- CP-element group 200: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1462_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1462_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1462_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1466_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1466_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1466_Sample/rr
      -- 
    ca_3372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1462_inst_ack_1, ack => convolution3D_CP_1767_elements(200)); -- 
    rr_3380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(200), ack => type_cast_1466_inst_req_0); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1466_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1466_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1466_Sample/ra
      -- 
    ra_3381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1466_inst_ack_0, ack => convolution3D_CP_1767_elements(201)); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	335 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1466_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1466_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1466_Update/ca
      -- 
    ca_3386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1466_inst_ack_1, ack => convolution3D_CP_1767_elements(202)); -- 
    -- CP-element group 203:  join  transition  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	186 
    -- CP-element group 203: 	170 
    -- CP-element group 203: 	182 
    -- CP-element group 203: 	174 
    -- CP-element group 203: 	178 
    -- CP-element group 203: 	190 
    -- CP-element group 203: 	194 
    -- CP-element group 203: 	198 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (9) 
      -- CP-element group 203: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Sample/ptr_deref_1474_Split/$entry
      -- CP-element group 203: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Sample/ptr_deref_1474_Split/$exit
      -- CP-element group 203: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Sample/ptr_deref_1474_Split/split_req
      -- CP-element group 203: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Sample/ptr_deref_1474_Split/split_ack
      -- CP-element group 203: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Sample/word_access_start/$entry
      -- CP-element group 203: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Sample/word_access_start/word_0/$entry
      -- CP-element group 203: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Sample/word_access_start/word_0/rr
      -- 
    rr_3424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(203), ack => ptr_deref_1474_store_0_req_0); -- 
    convolution3D_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(186) & convolution3D_CP_1767_elements(170) & convolution3D_CP_1767_elements(182) & convolution3D_CP_1767_elements(174) & convolution3D_CP_1767_elements(178) & convolution3D_CP_1767_elements(190) & convolution3D_CP_1767_elements(194) & convolution3D_CP_1767_elements(198) & convolution3D_CP_1767_elements(202);
      gj_convolution3D_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (5) 
      -- CP-element group 204: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Sample/word_access_start/$exit
      -- CP-element group 204: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Sample/word_access_start/word_0/$exit
      -- CP-element group 204: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Sample/word_access_start/word_0/ra
      -- 
    ra_3425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1474_store_0_ack_0, ack => convolution3D_CP_1767_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	335 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (5) 
      -- CP-element group 205: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Update/word_access_complete/$exit
      -- CP-element group 205: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Update/word_access_complete/word_0/$exit
      -- CP-element group 205: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Update/word_access_complete/word_0/ca
      -- 
    ca_3436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1474_store_0_ack_1, ack => convolution3D_CP_1767_elements(205)); -- 
    -- CP-element group 206:  branch  join  transition  place  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	167 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206: 	208 
    -- CP-element group 206:  members (10) 
      -- CP-element group 206: 	 branch_block_stmt_554/if_stmt_1488_eval_test/$entry
      -- CP-element group 206: 	 branch_block_stmt_554/if_stmt_1488__entry__
      -- CP-element group 206: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487__exit__
      -- CP-element group 206: 	 branch_block_stmt_554/if_stmt_1488_eval_test/$exit
      -- CP-element group 206: 	 branch_block_stmt_554/if_stmt_1488_eval_test/branch_req
      -- CP-element group 206: 	 branch_block_stmt_554/if_stmt_1488_if_link/$entry
      -- CP-element group 206: 	 branch_block_stmt_554/if_stmt_1488_else_link/$entry
      -- CP-element group 206: 	 branch_block_stmt_554/R_exitcond_1489_place
      -- CP-element group 206: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/$exit
      -- CP-element group 206: 	 branch_block_stmt_554/if_stmt_1488_dead_link/$entry
      -- 
    branch_req_3444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(206), ack => if_stmt_1488_branch_req_0); -- 
    convolution3D_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(167) & convolution3D_CP_1767_elements(205);
      gj_convolution3D_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	336 
    -- CP-element group 207: 	337 
    -- CP-element group 207:  members (24) 
      -- CP-element group 207: 	 branch_block_stmt_554/assign_stmt_1501_to_assign_stmt_1516__exit__
      -- CP-element group 207: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215
      -- CP-element group 207: 	 branch_block_stmt_554/assign_stmt_1501_to_assign_stmt_1516__entry__
      -- CP-element group 207: 	 branch_block_stmt_554/merge_stmt_1494__exit__
      -- CP-element group 207: 	 branch_block_stmt_554/if_stmt_1488_if_link/$exit
      -- CP-element group 207: 	 branch_block_stmt_554/if_stmt_1488_if_link/if_choice_transition
      -- CP-element group 207: 	 branch_block_stmt_554/assign_stmt_1501_to_assign_stmt_1516/$entry
      -- CP-element group 207: 	 branch_block_stmt_554/assign_stmt_1501_to_assign_stmt_1516/$exit
      -- CP-element group 207: 	 branch_block_stmt_554/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge
      -- CP-element group 207: 	 branch_block_stmt_554/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge_PhiReq/$entry
      -- CP-element group 207: 	 branch_block_stmt_554/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge_PhiReq/$exit
      -- CP-element group 207: 	 branch_block_stmt_554/merge_stmt_1494_PhiReqMerge
      -- CP-element group 207: 	 branch_block_stmt_554/merge_stmt_1494_PhiAck/$entry
      -- CP-element group 207: 	 branch_block_stmt_554/merge_stmt_1494_PhiAck/$exit
      -- CP-element group 207: 	 branch_block_stmt_554/merge_stmt_1494_PhiAck/dummy
      -- CP-element group 207: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/$entry
      -- CP-element group 207: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1519/$entry
      -- CP-element group 207: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/$entry
      -- CP-element group 207: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/$entry
      -- CP-element group 207: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/$entry
      -- CP-element group 207: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/Sample/rr
      -- CP-element group 207: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/Update/cr
      -- 
    if_choice_transition_3449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1488_branch_ack_1, ack => convolution3D_CP_1767_elements(207)); -- 
    rr_4425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(207), ack => type_cast_1522_inst_req_0); -- 
    cr_4430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(207), ack => type_cast_1522_inst_req_1); -- 
    -- CP-element group 208:  fork  transition  place  input  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	331 
    -- CP-element group 208: 	332 
    -- CP-element group 208:  members (12) 
      -- CP-element group 208: 	 branch_block_stmt_554/if_stmt_1488_else_link/$exit
      -- CP-element group 208: 	 branch_block_stmt_554/if_stmt_1488_else_link/else_choice_transition
      -- CP-element group 208: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163
      -- CP-element group 208: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/$entry
      -- CP-element group 208: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1325/$entry
      -- CP-element group 208: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_sources/$entry
      -- CP-element group 208: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_sources/type_cast_1331/$entry
      -- CP-element group 208: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_sources/type_cast_1331/SplitProtocol/$entry
      -- CP-element group 208: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_sources/type_cast_1331/SplitProtocol/Sample/$entry
      -- CP-element group 208: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_sources/type_cast_1331/SplitProtocol/Sample/rr
      -- CP-element group 208: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_sources/type_cast_1331/SplitProtocol/Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_sources/type_cast_1331/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1488_branch_ack_0, ack => convolution3D_CP_1767_elements(208)); -- 
    rr_4382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(208), ack => type_cast_1331_inst_req_0); -- 
    cr_4387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(208), ack => type_cast_1331_inst_req_1); -- 
    -- CP-element group 209:  transition  place  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	341 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	360 
    -- CP-element group 209:  members (5) 
      -- CP-element group 209: 	 branch_block_stmt_554/forx_xend215_ifx_xend227
      -- CP-element group 209: 	 branch_block_stmt_554/if_stmt_1539_if_link/if_choice_transition
      -- CP-element group 209: 	 branch_block_stmt_554/if_stmt_1539_if_link/$exit
      -- CP-element group 209: 	 branch_block_stmt_554/forx_xend215_ifx_xend227_PhiReq/$exit
      -- CP-element group 209: 	 branch_block_stmt_554/forx_xend215_ifx_xend227_PhiReq/$entry
      -- 
    if_choice_transition_3474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1539_branch_ack_1, ack => convolution3D_CP_1767_elements(209)); -- 
    -- CP-element group 210:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	341 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (18) 
      -- CP-element group 210: 	 branch_block_stmt_554/if_stmt_1539_else_link/else_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_554/assign_stmt_1551_to_assign_stmt_1561__entry__
      -- CP-element group 210: 	 branch_block_stmt_554/merge_stmt_1545__exit__
      -- CP-element group 210: 	 branch_block_stmt_554/if_stmt_1539_else_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_554/assign_stmt_1551_to_assign_stmt_1561/$entry
      -- CP-element group 210: 	 branch_block_stmt_554/forx_xend215_bbx_xnphx_xi340
      -- CP-element group 210: 	 branch_block_stmt_554/assign_stmt_1551_to_assign_stmt_1561/type_cast_1554_Update/cr
      -- CP-element group 210: 	 branch_block_stmt_554/assign_stmt_1551_to_assign_stmt_1561/type_cast_1554_Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_554/assign_stmt_1551_to_assign_stmt_1561/type_cast_1554_Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_554/assign_stmt_1551_to_assign_stmt_1561/type_cast_1554_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_554/assign_stmt_1551_to_assign_stmt_1561/type_cast_1554_update_start_
      -- CP-element group 210: 	 branch_block_stmt_554/assign_stmt_1551_to_assign_stmt_1561/type_cast_1554_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_554/forx_xend215_bbx_xnphx_xi340_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_554/forx_xend215_bbx_xnphx_xi340_PhiReq/$exit
      -- CP-element group 210: 	 branch_block_stmt_554/merge_stmt_1545_PhiReqMerge
      -- CP-element group 210: 	 branch_block_stmt_554/merge_stmt_1545_PhiAck/$entry
      -- CP-element group 210: 	 branch_block_stmt_554/merge_stmt_1545_PhiAck/$exit
      -- CP-element group 210: 	 branch_block_stmt_554/merge_stmt_1545_PhiAck/dummy
      -- 
    else_choice_transition_3478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1539_branch_ack_0, ack => convolution3D_CP_1767_elements(210)); -- 
    cr_3496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(210), ack => type_cast_1554_inst_req_1); -- 
    rr_3491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(210), ack => type_cast_1554_inst_req_0); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_554/assign_stmt_1551_to_assign_stmt_1561/type_cast_1554_Sample/ra
      -- CP-element group 211: 	 branch_block_stmt_554/assign_stmt_1551_to_assign_stmt_1561/type_cast_1554_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_554/assign_stmt_1551_to_assign_stmt_1561/type_cast_1554_sample_completed_
      -- 
    ra_3492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1554_inst_ack_0, ack => convolution3D_CP_1767_elements(211)); -- 
    -- CP-element group 212:  fork  transition  place  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	342 
    -- CP-element group 212: 	343 
    -- CP-element group 212:  members (11) 
      -- CP-element group 212: 	 branch_block_stmt_554/bbx_xnphx_xi340_forx_xbodyx_xi349
      -- CP-element group 212: 	 branch_block_stmt_554/assign_stmt_1551_to_assign_stmt_1561__exit__
      -- CP-element group 212: 	 branch_block_stmt_554/assign_stmt_1551_to_assign_stmt_1561/type_cast_1554_Update/ca
      -- CP-element group 212: 	 branch_block_stmt_554/assign_stmt_1551_to_assign_stmt_1561/type_cast_1554_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_554/assign_stmt_1551_to_assign_stmt_1561/type_cast_1554_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_554/assign_stmt_1551_to_assign_stmt_1561/$exit
      -- CP-element group 212: 	 branch_block_stmt_554/bbx_xnphx_xi340_forx_xbodyx_xi349_PhiReq/$entry
      -- CP-element group 212: 	 branch_block_stmt_554/bbx_xnphx_xi340_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/$entry
      -- CP-element group 212: 	 branch_block_stmt_554/bbx_xnphx_xi340_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/$entry
      -- CP-element group 212: 	 branch_block_stmt_554/bbx_xnphx_xi340_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/$entry
      -- CP-element group 212: 	 branch_block_stmt_554/bbx_xnphx_xi340_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_sources/$entry
      -- 
    ca_3497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1554_inst_ack_1, ack => convolution3D_CP_1767_elements(212)); -- 
    -- CP-element group 213:  transition  input  output  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	355 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213:  members (6) 
      -- CP-element group 213: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/RPIPE_maxpool_input_pipe_1592_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/RPIPE_maxpool_input_pipe_1592_update_start_
      -- CP-element group 213: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/RPIPE_maxpool_input_pipe_1592_Update/cr
      -- CP-element group 213: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/RPIPE_maxpool_input_pipe_1592_Update/$entry
      -- CP-element group 213: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/RPIPE_maxpool_input_pipe_1592_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/RPIPE_maxpool_input_pipe_1592_Sample/ra
      -- 
    ra_3509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1592_inst_ack_0, ack => convolution3D_CP_1767_elements(213)); -- 
    cr_3513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(213), ack => RPIPE_maxpool_input_pipe_1592_inst_req_1); -- 
    -- CP-element group 214:  transition  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	213 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (6) 
      -- CP-element group 214: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1596_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/RPIPE_maxpool_input_pipe_1592_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/RPIPE_maxpool_input_pipe_1592_Update/ca
      -- CP-element group 214: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/RPIPE_maxpool_input_pipe_1592_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1596_Sample/rr
      -- CP-element group 214: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1596_Sample/$entry
      -- 
    ca_3514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1592_inst_ack_1, ack => convolution3D_CP_1767_elements(214)); -- 
    rr_3522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(214), ack => type_cast_1596_inst_req_0); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1596_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1596_Sample/ra
      -- CP-element group 215: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1596_Sample/$exit
      -- 
    ra_3523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1596_inst_ack_0, ack => convolution3D_CP_1767_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	355 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	219 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1596_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1596_Update/ca
      -- CP-element group 216: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1596_Update/$exit
      -- 
    ca_3528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1596_inst_ack_1, ack => convolution3D_CP_1767_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	355 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1611_Sample/ra
      -- CP-element group 217: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1611_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1611_sample_completed_
      -- 
    ra_3537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1611_inst_ack_0, ack => convolution3D_CP_1767_elements(217)); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	355 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1611_Update/ca
      -- CP-element group 218: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1611_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1611_update_completed_
      -- 
    ca_3542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1611_inst_ack_1, ack => convolution3D_CP_1767_elements(218)); -- 
    -- CP-element group 219:  branch  join  transition  place  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: 	216 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (10) 
      -- CP-element group 219: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617__exit__
      -- CP-element group 219: 	 branch_block_stmt_554/if_stmt_1618__entry__
      -- CP-element group 219: 	 branch_block_stmt_554/R_cmpx_xi348_1619_place
      -- CP-element group 219: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/$exit
      -- CP-element group 219: 	 branch_block_stmt_554/if_stmt_1618_else_link/$entry
      -- CP-element group 219: 	 branch_block_stmt_554/if_stmt_1618_if_link/$entry
      -- CP-element group 219: 	 branch_block_stmt_554/if_stmt_1618_eval_test/branch_req
      -- CP-element group 219: 	 branch_block_stmt_554/if_stmt_1618_eval_test/$exit
      -- CP-element group 219: 	 branch_block_stmt_554/if_stmt_1618_eval_test/$entry
      -- CP-element group 219: 	 branch_block_stmt_554/if_stmt_1618_dead_link/$entry
      -- 
    branch_req_3550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(219), ack => if_stmt_1618_branch_req_0); -- 
    convolution3D_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(218) & convolution3D_CP_1767_elements(216);
      gj_convolution3D_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  fork  transition  place  input  output  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	345 
    -- CP-element group 220: 	346 
    -- CP-element group 220: 	348 
    -- CP-element group 220: 	349 
    -- CP-element group 220:  members (20) 
      -- CP-element group 220: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349
      -- CP-element group 220: 	 branch_block_stmt_554/if_stmt_1618_if_link/if_choice_transition
      -- CP-element group 220: 	 branch_block_stmt_554/if_stmt_1618_if_link/$exit
      -- CP-element group 220: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1570/SplitProtocol/$entry
      -- CP-element group 220: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1570/SplitProtocol/Sample/$entry
      -- CP-element group 220: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_sources/type_cast_1577/SplitProtocol/Sample/$entry
      -- CP-element group 220: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1570/$entry
      -- CP-element group 220: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/$entry
      -- CP-element group 220: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_sources/type_cast_1577/SplitProtocol/$entry
      -- CP-element group 220: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_sources/type_cast_1577/$entry
      -- CP-element group 220: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_sources/$entry
      -- CP-element group 220: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/$entry
      -- CP-element group 220: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/$entry
      -- CP-element group 220: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1570/SplitProtocol/Update/cr
      -- CP-element group 220: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1570/SplitProtocol/Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1570/SplitProtocol/Sample/rr
      -- CP-element group 220: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/$entry
      -- CP-element group 220: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_sources/type_cast_1577/SplitProtocol/Update/cr
      -- CP-element group 220: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_sources/type_cast_1577/SplitProtocol/Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_sources/type_cast_1577/SplitProtocol/Sample/rr
      -- 
    if_choice_transition_3555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1618_branch_ack_1, ack => convolution3D_CP_1767_elements(220)); -- 
    cr_4503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(220), ack => type_cast_1570_inst_req_1); -- 
    rr_4498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(220), ack => type_cast_1570_inst_req_0); -- 
    cr_4526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(220), ack => type_cast_1577_inst_req_1); -- 
    rr_4521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(220), ack => type_cast_1577_inst_req_0); -- 
    -- CP-element group 221:  fork  transition  place  input  output  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	356 
    -- CP-element group 221: 	357 
    -- CP-element group 221:  members (12) 
      -- CP-element group 221: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357
      -- CP-element group 221: 	 branch_block_stmt_554/if_stmt_1618_else_link/else_choice_transition
      -- CP-element group 221: 	 branch_block_stmt_554/if_stmt_1618_else_link/$exit
      -- CP-element group 221: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1628/SplitProtocol/$entry
      -- CP-element group 221: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1628/SplitProtocol/Sample/$entry
      -- CP-element group 221: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1628/$entry
      -- CP-element group 221: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/$entry
      -- CP-element group 221: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/phi_stmt_1625/$entry
      -- CP-element group 221: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1628/SplitProtocol/Update/cr
      -- CP-element group 221: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1628/SplitProtocol/Update/$entry
      -- CP-element group 221: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1628/SplitProtocol/Sample/rr
      -- 
    else_choice_transition_3559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1618_branch_ack_0, ack => convolution3D_CP_1767_elements(221)); -- 
    cr_4562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(221), ack => type_cast_1628_inst_req_1); -- 
    rr_4557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(221), ack => type_cast_1628_inst_req_0); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	359 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	228 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_final_index_sum_regn_sample_complete
      -- CP-element group 222: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_final_index_sum_regn_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_final_index_sum_regn_Sample/ack
      -- 
    ack_3590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1657_index_offset_ack_0, ack => convolution3D_CP_1767_elements(222)); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	359 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (11) 
      -- CP-element group 223: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_base_plus_offset/sum_rename_ack
      -- CP-element group 223: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/addr_of_1658_request/$entry
      -- CP-element group 223: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_base_plus_offset/sum_rename_req
      -- CP-element group 223: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_base_plus_offset/$exit
      -- CP-element group 223: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_base_plus_offset/$entry
      -- CP-element group 223: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_offset_calculated
      -- CP-element group 223: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_final_index_sum_regn_Update/ack
      -- CP-element group 223: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_root_address_calculated
      -- CP-element group 223: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_final_index_sum_regn_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/addr_of_1658_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/addr_of_1658_request/req
      -- 
    ack_3595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1657_index_offset_ack_1, ack => convolution3D_CP_1767_elements(223)); -- 
    req_3604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(223), ack => addr_of_1658_final_reg_req_0); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/addr_of_1658_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/addr_of_1658_request/ack
      -- CP-element group 224: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/addr_of_1658_request/$exit
      -- 
    ack_3605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1658_final_reg_ack_0, ack => convolution3D_CP_1767_elements(224)); -- 
    -- CP-element group 225:  join  fork  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	359 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (28) 
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Sample/word_access_start/word_0/rr
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Sample/word_access_start/word_0/$entry
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Sample/word_access_start/$entry
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/addr_of_1658_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Sample/ptr_deref_1661_Split/split_ack
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Sample/ptr_deref_1661_Split/split_req
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Sample/ptr_deref_1661_Split/$exit
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Sample/ptr_deref_1661_Split/$entry
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_word_addrgen/root_register_ack
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_word_addrgen/root_register_req
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_word_addrgen/$exit
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_word_addrgen/$entry
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_base_plus_offset/$entry
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_base_addr_resize/base_resize_ack
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_base_addr_resize/base_resize_req
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_base_addr_resize/$exit
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_base_addr_resize/$entry
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_base_address_resized
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_word_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_base_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/addr_of_1658_complete/ack
      -- CP-element group 225: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/addr_of_1658_complete/$exit
      -- 
    ack_3610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1658_final_reg_ack_1, ack => convolution3D_CP_1767_elements(225)); -- 
    rr_3648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(225), ack => ptr_deref_1661_store_0_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (5) 
      -- CP-element group 226: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Sample/word_access_start/word_0/ra
      -- CP-element group 226: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Sample/word_access_start/word_0/$exit
      -- CP-element group 226: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Sample/word_access_start/$exit
      -- CP-element group 226: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_sample_completed_
      -- 
    ra_3649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1661_store_0_ack_0, ack => convolution3D_CP_1767_elements(226)); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	359 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Update/word_access_complete/word_0/ca
      -- CP-element group 227: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Update/word_access_complete/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Update/word_access_complete/$exit
      -- CP-element group 227: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_update_completed_
      -- 
    ca_3660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1661_store_0_ack_1, ack => convolution3D_CP_1767_elements(227)); -- 
    -- CP-element group 228:  join  transition  place  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	222 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	360 
    -- CP-element group 228:  members (5) 
      -- CP-element group 228: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663__exit__
      -- CP-element group 228: 	 branch_block_stmt_554/getRemainingElementsx_xexit357_ifx_xend227
      -- CP-element group 228: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/$exit
      -- CP-element group 228: 	 branch_block_stmt_554/getRemainingElementsx_xexit357_ifx_xend227_PhiReq/$exit
      -- CP-element group 228: 	 branch_block_stmt_554/getRemainingElementsx_xexit357_ifx_xend227_PhiReq/$entry
      -- 
    convolution3D_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(222) & convolution3D_CP_1767_elements(227);
      gj_convolution3D_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  transition  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	360 
    -- CP-element group 229: successors 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_554/call_stmt_1668/call_stmt_1668_Sample/$exit
      -- CP-element group 229: 	 branch_block_stmt_554/call_stmt_1668/call_stmt_1668_Sample/cra
      -- CP-element group 229: 	 branch_block_stmt_554/call_stmt_1668/call_stmt_1668_sample_completed_
      -- 
    cra_3672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1668_call_ack_0, ack => convolution3D_CP_1767_elements(229)); -- 
    -- CP-element group 230:  fork  transition  place  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	360 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	237 
    -- CP-element group 230: 	238 
    -- CP-element group 230: 	235 
    -- CP-element group 230: 	236 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (22) 
      -- CP-element group 230: 	 branch_block_stmt_554/call_stmt_1668__exit__
      -- CP-element group 230: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707__entry__
      -- CP-element group 230: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1701_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_554/call_stmt_1668/call_stmt_1668_update_completed_
      -- CP-element group 230: 	 branch_block_stmt_554/call_stmt_1668/$exit
      -- CP-element group 230: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1691_Update/cr
      -- CP-element group 230: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1691_Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1691_Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1691_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1691_update_start_
      -- CP-element group 230: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1691_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/$entry
      -- CP-element group 230: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1670_Sample/req
      -- CP-element group 230: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1670_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1670_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1701_Update/cr
      -- CP-element group 230: 	 branch_block_stmt_554/call_stmt_1668/call_stmt_1668_Update/cca
      -- CP-element group 230: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1701_Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1701_Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1701_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_554/call_stmt_1668/call_stmt_1668_Update/$exit
      -- CP-element group 230: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1701_update_start_
      -- 
    cca_3677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1668_call_ack_1, ack => convolution3D_CP_1767_elements(230)); -- 
    cr_3721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(230), ack => type_cast_1691_inst_req_1); -- 
    rr_3716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(230), ack => type_cast_1691_inst_req_0); -- 
    req_3688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(230), ack => WPIPE_maxpool_output_pipe_1670_inst_req_0); -- 
    cr_3735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(230), ack => type_cast_1701_inst_req_1); -- 
    rr_3730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(230), ack => type_cast_1701_inst_req_0); -- 
    -- CP-element group 231:  transition  input  output  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (6) 
      -- CP-element group 231: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1670_Update/req
      -- CP-element group 231: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1670_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1670_Sample/ack
      -- CP-element group 231: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1670_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1670_update_start_
      -- CP-element group 231: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1670_sample_completed_
      -- 
    ack_3689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1670_inst_ack_0, ack => convolution3D_CP_1767_elements(231)); -- 
    req_3693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(231), ack => WPIPE_maxpool_output_pipe_1670_inst_req_1); -- 
    -- CP-element group 232:  transition  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	233 
    -- CP-element group 232:  members (6) 
      -- CP-element group 232: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1674_Sample/req
      -- CP-element group 232: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1674_Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1674_sample_start_
      -- CP-element group 232: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1670_Update/ack
      -- CP-element group 232: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1670_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1670_update_completed_
      -- 
    ack_3694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1670_inst_ack_1, ack => convolution3D_CP_1767_elements(232)); -- 
    req_3702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(232), ack => WPIPE_maxpool_output_pipe_1674_inst_req_0); -- 
    -- CP-element group 233:  transition  input  output  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	232 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	234 
    -- CP-element group 233:  members (6) 
      -- CP-element group 233: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1674_Update/req
      -- CP-element group 233: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1674_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1674_Sample/ack
      -- CP-element group 233: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1674_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1674_update_start_
      -- CP-element group 233: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1674_sample_completed_
      -- 
    ack_3703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1674_inst_ack_0, ack => convolution3D_CP_1767_elements(233)); -- 
    req_3707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(233), ack => WPIPE_maxpool_output_pipe_1674_inst_req_1); -- 
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	233 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	239 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1674_Update/ack
      -- CP-element group 234: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1674_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/WPIPE_maxpool_output_pipe_1674_update_completed_
      -- 
    ack_3708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1674_inst_ack_1, ack => convolution3D_CP_1767_elements(234)); -- 
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	230 
    -- CP-element group 235: successors 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1691_Sample/ra
      -- CP-element group 235: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1691_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1691_sample_completed_
      -- 
    ra_3717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1691_inst_ack_0, ack => convolution3D_CP_1767_elements(235)); -- 
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	230 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	239 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1691_Update/ca
      -- CP-element group 236: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1691_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1691_update_completed_
      -- 
    ca_3722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1691_inst_ack_1, ack => convolution3D_CP_1767_elements(236)); -- 
    -- CP-element group 237:  transition  input  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	230 
    -- CP-element group 237: successors 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1701_Sample/ra
      -- CP-element group 237: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1701_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1701_sample_completed_
      -- 
    ra_3731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1701_inst_ack_0, ack => convolution3D_CP_1767_elements(237)); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	230 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1701_Update/ca
      -- CP-element group 238: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1701_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/type_cast_1701_update_completed_
      -- 
    ca_3736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1701_inst_ack_1, ack => convolution3D_CP_1767_elements(238)); -- 
    -- CP-element group 239:  join  transition  place  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: 	234 
    -- CP-element group 239: 	236 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	361 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_554/ifx_xend227_whilex_xbody
      -- CP-element group 239: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707__exit__
      -- CP-element group 239: 	 branch_block_stmt_554/assign_stmt_1673_to_assign_stmt_1707/$exit
      -- CP-element group 239: 	 branch_block_stmt_554/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_sources/$entry
      -- CP-element group 239: 	 branch_block_stmt_554/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1710/$entry
      -- CP-element group 239: 	 branch_block_stmt_554/ifx_xend227_whilex_xbody_PhiReq/$entry
      -- 
    convolution3D_cp_element_group_239: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_239"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(238) & convolution3D_CP_1767_elements(234) & convolution3D_CP_1767_elements(236);
      gj_convolution3D_cp_element_group_239 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(239), clk => clk, reset => reset); --
    end block;
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	366 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1723_Sample/ack
      -- CP-element group 240: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1723_Update/$entry
      -- CP-element group 240: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1723_Update/req
      -- CP-element group 240: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1723_Sample/$exit
      -- CP-element group 240: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1723_update_start_
      -- CP-element group 240: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1723_sample_completed_
      -- 
    ack_3748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1723_inst_ack_0, ack => convolution3D_CP_1767_elements(240)); -- 
    req_3752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(240), ack => WPIPE_num_out_pipe_1723_inst_req_1); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1723_Update/ack
      -- CP-element group 241: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1723_Update/$exit
      -- CP-element group 241: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1726_Sample/req
      -- CP-element group 241: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1726_Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1723_update_completed_
      -- CP-element group 241: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1726_sample_start_
      -- 
    ack_3753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1723_inst_ack_1, ack => convolution3D_CP_1767_elements(241)); -- 
    req_3761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(241), ack => WPIPE_num_out_pipe_1726_inst_req_0); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1726_Sample/ack
      -- CP-element group 242: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1726_Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1726_Sample/$exit
      -- CP-element group 242: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1726_update_start_
      -- CP-element group 242: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1726_sample_completed_
      -- CP-element group 242: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1726_Update/req
      -- 
    ack_3762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1726_inst_ack_0, ack => convolution3D_CP_1767_elements(242)); -- 
    req_3766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(242), ack => WPIPE_num_out_pipe_1726_inst_req_1); -- 
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	248 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1726_update_completed_
      -- CP-element group 243: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1726_Update/ack
      -- CP-element group 243: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1726_Update/$exit
      -- 
    ack_3767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1726_inst_ack_1, ack => convolution3D_CP_1767_elements(243)); -- 
    -- CP-element group 244:  transition  input  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	366 
    -- CP-element group 244: successors 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1737_Sample/cra
      -- CP-element group 244: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1737_Sample/$exit
      -- CP-element group 244: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1737_sample_completed_
      -- 
    cra_3776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1737_call_ack_0, ack => convolution3D_CP_1767_elements(244)); -- 
    -- CP-element group 245:  transition  input  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	366 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	248 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1737_Update/cca
      -- CP-element group 245: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1737_Update/$exit
      -- CP-element group 245: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1737_update_completed_
      -- 
    cca_3781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1737_call_ack_1, ack => convolution3D_CP_1767_elements(245)); -- 
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	366 
    -- CP-element group 246: successors 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1741_Sample/cra
      -- CP-element group 246: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1741_Sample/$exit
      -- CP-element group 246: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1741_sample_completed_
      -- 
    cra_3790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1741_call_ack_0, ack => convolution3D_CP_1767_elements(246)); -- 
    -- CP-element group 247:  transition  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	366 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1741_Update/cca
      -- CP-element group 247: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1741_Update/$exit
      -- CP-element group 247: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1741_update_completed_
      -- 
    cca_3795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1741_call_ack_1, ack => convolution3D_CP_1767_elements(247)); -- 
    -- CP-element group 248:  branch  join  transition  place  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	245 
    -- CP-element group 248: 	247 
    -- CP-element group 248: 	243 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248: 	250 
    -- CP-element group 248:  members (10) 
      -- CP-element group 248: 	 branch_block_stmt_554/R_exitcond5_1754_place
      -- CP-element group 248: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752__exit__
      -- CP-element group 248: 	 branch_block_stmt_554/if_stmt_1753__entry__
      -- CP-element group 248: 	 branch_block_stmt_554/if_stmt_1753_eval_test/branch_req
      -- CP-element group 248: 	 branch_block_stmt_554/if_stmt_1753_if_link/$entry
      -- CP-element group 248: 	 branch_block_stmt_554/if_stmt_1753_eval_test/$exit
      -- CP-element group 248: 	 branch_block_stmt_554/if_stmt_1753_eval_test/$entry
      -- CP-element group 248: 	 branch_block_stmt_554/if_stmt_1753_dead_link/$entry
      -- CP-element group 248: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/$exit
      -- CP-element group 248: 	 branch_block_stmt_554/if_stmt_1753_else_link/$entry
      -- 
    branch_req_3803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(248), ack => if_stmt_1753_branch_req_0); -- 
    convolution3D_cp_element_group_248: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_248"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(245) & convolution3D_CP_1767_elements(247) & convolution3D_CP_1767_elements(243);
      gj_convolution3D_cp_element_group_248 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(248), clk => clk, reset => reset); --
    end block;
    -- CP-element group 249:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	253 
    -- CP-element group 249: 	251 
    -- CP-element group 249: 	252 
    -- CP-element group 249:  members (21) 
      -- CP-element group 249: 	 branch_block_stmt_554/whilex_xbody_whilex_xend
      -- CP-element group 249: 	 branch_block_stmt_554/merge_stmt_1759_PhiReqMerge
      -- CP-element group 249: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767__entry__
      -- CP-element group 249: 	 branch_block_stmt_554/merge_stmt_1759__exit__
      -- CP-element group 249: 	 branch_block_stmt_554/if_stmt_1753_if_link/$exit
      -- CP-element group 249: 	 branch_block_stmt_554/if_stmt_1753_if_link/if_choice_transition
      -- CP-element group 249: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/RPIPE_input_done_pipe_1766_Sample/rr
      -- CP-element group 249: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/RPIPE_input_done_pipe_1766_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/type_cast_1763_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/$entry
      -- CP-element group 249: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/RPIPE_input_done_pipe_1766_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/type_cast_1763_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/type_cast_1763_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/type_cast_1763_Sample/rr
      -- CP-element group 249: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/type_cast_1763_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/type_cast_1763_update_start_
      -- CP-element group 249: 	 branch_block_stmt_554/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 249: 	 branch_block_stmt_554/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 249: 	 branch_block_stmt_554/merge_stmt_1759_PhiAck/$entry
      -- CP-element group 249: 	 branch_block_stmt_554/merge_stmt_1759_PhiAck/$exit
      -- CP-element group 249: 	 branch_block_stmt_554/merge_stmt_1759_PhiAck/dummy
      -- 
    if_choice_transition_3808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1753_branch_ack_1, ack => convolution3D_CP_1767_elements(249)); -- 
    rr_3839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(249), ack => RPIPE_input_done_pipe_1766_inst_req_0); -- 
    cr_3830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(249), ack => type_cast_1763_inst_req_1); -- 
    rr_3825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(249), ack => type_cast_1763_inst_req_0); -- 
    -- CP-element group 250:  fork  transition  place  input  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	248 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	362 
    -- CP-element group 250: 	363 
    -- CP-element group 250:  members (12) 
      -- CP-element group 250: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody
      -- CP-element group 250: 	 branch_block_stmt_554/if_stmt_1753_else_link/else_choice_transition
      -- CP-element group 250: 	 branch_block_stmt_554/if_stmt_1753_else_link/$exit
      -- CP-element group 250: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_sources/type_cast_1713/SplitProtocol/Update/cr
      -- CP-element group 250: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_sources/type_cast_1713/SplitProtocol/Update/$entry
      -- CP-element group 250: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_sources/type_cast_1713/SplitProtocol/Sample/rr
      -- CP-element group 250: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_sources/type_cast_1713/SplitProtocol/Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_sources/type_cast_1713/SplitProtocol/$entry
      -- CP-element group 250: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_sources/type_cast_1713/$entry
      -- CP-element group 250: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_sources/$entry
      -- CP-element group 250: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1710/$entry
      -- CP-element group 250: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/$entry
      -- 
    else_choice_transition_3812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1753_branch_ack_0, ack => convolution3D_CP_1767_elements(250)); -- 
    cr_4615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(250), ack => type_cast_1713_inst_req_1); -- 
    rr_4610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(250), ack => type_cast_1713_inst_req_0); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: successors 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/type_cast_1763_Sample/ra
      -- CP-element group 251: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/type_cast_1763_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/type_cast_1763_sample_completed_
      -- 
    ra_3826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1763_inst_ack_0, ack => convolution3D_CP_1767_elements(251)); -- 
    -- CP-element group 252:  transition  input  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	249 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	255 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/type_cast_1763_Update/ca
      -- CP-element group 252: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/type_cast_1763_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/type_cast_1763_update_completed_
      -- 
    ca_3831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1763_inst_ack_1, ack => convolution3D_CP_1767_elements(252)); -- 
    -- CP-element group 253:  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	249 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/RPIPE_input_done_pipe_1766_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/RPIPE_input_done_pipe_1766_update_start_
      -- CP-element group 253: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/RPIPE_input_done_pipe_1766_sample_completed_
      -- CP-element group 253: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/RPIPE_input_done_pipe_1766_Update/cr
      -- CP-element group 253: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/RPIPE_input_done_pipe_1766_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/RPIPE_input_done_pipe_1766_Sample/ra
      -- 
    ra_3840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_1766_inst_ack_0, ack => convolution3D_CP_1767_elements(253)); -- 
    cr_3844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(253), ack => RPIPE_input_done_pipe_1766_inst_req_1); -- 
    -- CP-element group 254:  transition  input  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/RPIPE_input_done_pipe_1766_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/RPIPE_input_done_pipe_1766_Update/ca
      -- CP-element group 254: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/RPIPE_input_done_pipe_1766_Update/$exit
      -- 
    ca_3845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_1766_inst_ack_1, ack => convolution3D_CP_1767_elements(254)); -- 
    -- CP-element group 255:  join  fork  transition  place  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: 	252 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	275 
    -- CP-element group 255: 	273 
    -- CP-element group 255: 	269 
    -- CP-element group 255: 	271 
    -- CP-element group 255: 	261 
    -- CP-element group 255: 	263 
    -- CP-element group 255: 	265 
    -- CP-element group 255: 	267 
    -- CP-element group 255: 	256 
    -- CP-element group 255: 	257 
    -- CP-element group 255: 	259 
    -- CP-element group 255:  members (37) 
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878__entry__
      -- CP-element group 255: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767__exit__
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/call_stmt_1770_Update/ccr
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/call_stmt_1770_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1783_update_start_
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/call_stmt_1770_Sample/crr
      -- CP-element group 255: 	 branch_block_stmt_554/assign_stmt_1764_to_assign_stmt_1767/$exit
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/call_stmt_1770_Sample/$entry
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1774_Update/cr
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/call_stmt_1770_update_start_
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1774_update_start_
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/call_stmt_1770_sample_start_
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/$entry
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1774_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1783_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1783_Update/cr
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1793_update_start_
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1793_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1793_Update/cr
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1803_update_start_
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1803_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1803_Update/cr
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1813_update_start_
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1813_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1813_Update/cr
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1823_update_start_
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1823_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1823_Update/cr
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1833_update_start_
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1833_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1833_Update/cr
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1843_update_start_
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1843_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1843_Update/cr
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1853_update_start_
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1853_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1853_Update/cr
      -- 
    ccr_3861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(255), ack => call_stmt_1770_call_req_1); -- 
    crr_3856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(255), ack => call_stmt_1770_call_req_0); -- 
    cr_3875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(255), ack => type_cast_1774_inst_req_1); -- 
    cr_3889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(255), ack => type_cast_1783_inst_req_1); -- 
    cr_3903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(255), ack => type_cast_1793_inst_req_1); -- 
    cr_3917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(255), ack => type_cast_1803_inst_req_1); -- 
    cr_3931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(255), ack => type_cast_1813_inst_req_1); -- 
    cr_3945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(255), ack => type_cast_1823_inst_req_1); -- 
    cr_3959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(255), ack => type_cast_1833_inst_req_1); -- 
    cr_3973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(255), ack => type_cast_1843_inst_req_1); -- 
    cr_3987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(255), ack => type_cast_1853_inst_req_1); -- 
    convolution3D_cp_element_group_255: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_255"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(254) & convolution3D_CP_1767_elements(252);
      gj_convolution3D_cp_element_group_255 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(255), clk => clk, reset => reset); --
    end block;
    -- CP-element group 256:  transition  input  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/call_stmt_1770_Sample/cra
      -- CP-element group 256: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/call_stmt_1770_Sample/$exit
      -- CP-element group 256: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/call_stmt_1770_sample_completed_
      -- 
    cra_3857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1770_call_ack_0, ack => convolution3D_CP_1767_elements(256)); -- 
    -- CP-element group 257:  transition  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	255 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (6) 
      -- CP-element group 257: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1774_sample_start_
      -- CP-element group 257: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1774_Sample/rr
      -- CP-element group 257: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/call_stmt_1770_Update/cca
      -- CP-element group 257: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/call_stmt_1770_Update/$exit
      -- CP-element group 257: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1774_Sample/$entry
      -- CP-element group 257: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/call_stmt_1770_update_completed_
      -- 
    cca_3862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1770_call_ack_1, ack => convolution3D_CP_1767_elements(257)); -- 
    rr_3870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(257), ack => type_cast_1774_inst_req_0); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1774_Sample/$exit
      -- CP-element group 258: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1774_Sample/ra
      -- CP-element group 258: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1774_sample_completed_
      -- 
    ra_3871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1774_inst_ack_0, ack => convolution3D_CP_1767_elements(258)); -- 
    -- CP-element group 259:  fork  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	255 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	274 
    -- CP-element group 259: 	272 
    -- CP-element group 259: 	268 
    -- CP-element group 259: 	270 
    -- CP-element group 259: 	260 
    -- CP-element group 259: 	262 
    -- CP-element group 259: 	264 
    -- CP-element group 259: 	266 
    -- CP-element group 259:  members (27) 
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1774_Update/ca
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1783_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1783_Sample/rr
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1783_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1774_update_completed_
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1774_Update/$exit
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1793_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1793_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1793_Sample/rr
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1803_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1803_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1803_Sample/rr
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1813_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1813_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1813_Sample/rr
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1823_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1823_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1823_Sample/rr
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1833_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1833_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1833_Sample/rr
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1843_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1843_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1843_Sample/rr
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1853_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1853_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1853_Sample/rr
      -- 
    ca_3876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1774_inst_ack_1, ack => convolution3D_CP_1767_elements(259)); -- 
    rr_3968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(259), ack => type_cast_1843_inst_req_0); -- 
    rr_3982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(259), ack => type_cast_1853_inst_req_0); -- 
    rr_3954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(259), ack => type_cast_1833_inst_req_0); -- 
    rr_3884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(259), ack => type_cast_1783_inst_req_0); -- 
    rr_3898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(259), ack => type_cast_1793_inst_req_0); -- 
    rr_3912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(259), ack => type_cast_1803_inst_req_0); -- 
    rr_3926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(259), ack => type_cast_1813_inst_req_0); -- 
    rr_3940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(259), ack => type_cast_1823_inst_req_0); -- 
    -- CP-element group 260:  transition  input  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1783_sample_completed_
      -- CP-element group 260: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1783_Sample/ra
      -- CP-element group 260: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1783_Sample/$exit
      -- 
    ra_3885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1783_inst_ack_0, ack => convolution3D_CP_1767_elements(260)); -- 
    -- CP-element group 261:  transition  input  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	255 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	296 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1783_update_completed_
      -- CP-element group 261: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1783_Update/$exit
      -- CP-element group 261: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1783_Update/ca
      -- 
    ca_3890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1783_inst_ack_1, ack => convolution3D_CP_1767_elements(261)); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	259 
    -- CP-element group 262: successors 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1793_sample_completed_
      -- CP-element group 262: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1793_Sample/$exit
      -- CP-element group 262: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1793_Sample/ra
      -- 
    ra_3899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1793_inst_ack_0, ack => convolution3D_CP_1767_elements(262)); -- 
    -- CP-element group 263:  transition  input  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	255 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	293 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1793_update_completed_
      -- CP-element group 263: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1793_Update/$exit
      -- CP-element group 263: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1793_Update/ca
      -- 
    ca_3904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1793_inst_ack_1, ack => convolution3D_CP_1767_elements(263)); -- 
    -- CP-element group 264:  transition  input  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	259 
    -- CP-element group 264: successors 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1803_sample_completed_
      -- CP-element group 264: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1803_Sample/$exit
      -- CP-element group 264: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1803_Sample/ra
      -- 
    ra_3913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1803_inst_ack_0, ack => convolution3D_CP_1767_elements(264)); -- 
    -- CP-element group 265:  transition  input  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	255 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	290 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1803_update_completed_
      -- CP-element group 265: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1803_Update/$exit
      -- CP-element group 265: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1803_Update/ca
      -- 
    ca_3918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1803_inst_ack_1, ack => convolution3D_CP_1767_elements(265)); -- 
    -- CP-element group 266:  transition  input  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	259 
    -- CP-element group 266: successors 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1813_sample_completed_
      -- CP-element group 266: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1813_Sample/$exit
      -- CP-element group 266: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1813_Sample/ra
      -- 
    ra_3927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1813_inst_ack_0, ack => convolution3D_CP_1767_elements(266)); -- 
    -- CP-element group 267:  transition  input  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	255 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	287 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1813_update_completed_
      -- CP-element group 267: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1813_Update/$exit
      -- CP-element group 267: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1813_Update/ca
      -- 
    ca_3932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1813_inst_ack_1, ack => convolution3D_CP_1767_elements(267)); -- 
    -- CP-element group 268:  transition  input  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	259 
    -- CP-element group 268: successors 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1823_sample_completed_
      -- CP-element group 268: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1823_Sample/$exit
      -- CP-element group 268: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1823_Sample/ra
      -- 
    ra_3941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1823_inst_ack_0, ack => convolution3D_CP_1767_elements(268)); -- 
    -- CP-element group 269:  transition  input  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	255 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	284 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1823_update_completed_
      -- CP-element group 269: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1823_Update/$exit
      -- CP-element group 269: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1823_Update/ca
      -- 
    ca_3946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1823_inst_ack_1, ack => convolution3D_CP_1767_elements(269)); -- 
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	259 
    -- CP-element group 270: successors 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1833_sample_completed_
      -- CP-element group 270: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1833_Sample/$exit
      -- CP-element group 270: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1833_Sample/ra
      -- 
    ra_3955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1833_inst_ack_0, ack => convolution3D_CP_1767_elements(270)); -- 
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	255 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	281 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1833_update_completed_
      -- CP-element group 271: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1833_Update/$exit
      -- CP-element group 271: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1833_Update/ca
      -- 
    ca_3960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1833_inst_ack_1, ack => convolution3D_CP_1767_elements(271)); -- 
    -- CP-element group 272:  transition  input  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	259 
    -- CP-element group 272: successors 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1843_sample_completed_
      -- CP-element group 272: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1843_Sample/$exit
      -- CP-element group 272: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1843_Sample/ra
      -- 
    ra_3969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1843_inst_ack_0, ack => convolution3D_CP_1767_elements(272)); -- 
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	255 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	278 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1843_update_completed_
      -- CP-element group 273: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1843_Update/$exit
      -- CP-element group 273: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1843_Update/ca
      -- 
    ca_3974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1843_inst_ack_1, ack => convolution3D_CP_1767_elements(273)); -- 
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	259 
    -- CP-element group 274: successors 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1853_sample_completed_
      -- CP-element group 274: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1853_Sample/$exit
      -- CP-element group 274: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1853_Sample/ra
      -- 
    ra_3983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1853_inst_ack_0, ack => convolution3D_CP_1767_elements(274)); -- 
    -- CP-element group 275:  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	255 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1853_update_completed_
      -- CP-element group 275: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1853_Update/$exit
      -- CP-element group 275: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/type_cast_1853_Update/ca
      -- CP-element group 275: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1855_sample_start_
      -- CP-element group 275: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1855_Sample/$entry
      -- CP-element group 275: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1855_Sample/req
      -- 
    ca_3988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1853_inst_ack_1, ack => convolution3D_CP_1767_elements(275)); -- 
    req_3996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(275), ack => WPIPE_maxpool_output_pipe_1855_inst_req_0); -- 
    -- CP-element group 276:  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1855_sample_completed_
      -- CP-element group 276: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1855_update_start_
      -- CP-element group 276: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1855_Sample/$exit
      -- CP-element group 276: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1855_Sample/ack
      -- CP-element group 276: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1855_Update/$entry
      -- CP-element group 276: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1855_Update/req
      -- 
    ack_3997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1855_inst_ack_0, ack => convolution3D_CP_1767_elements(276)); -- 
    req_4001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(276), ack => WPIPE_maxpool_output_pipe_1855_inst_req_1); -- 
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1855_update_completed_
      -- CP-element group 277: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1855_Update/$exit
      -- CP-element group 277: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1855_Update/ack
      -- 
    ack_4002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1855_inst_ack_1, ack => convolution3D_CP_1767_elements(277)); -- 
    -- CP-element group 278:  join  transition  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: 	273 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1858_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1858_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1858_Sample/req
      -- 
    req_4010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(278), ack => WPIPE_maxpool_output_pipe_1858_inst_req_0); -- 
    convolution3D_cp_element_group_278: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_278"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(277) & convolution3D_CP_1767_elements(273);
      gj_convolution3D_cp_element_group_278 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(278), clk => clk, reset => reset); --
    end block;
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1858_sample_completed_
      -- CP-element group 279: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1858_update_start_
      -- CP-element group 279: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1858_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1858_Sample/ack
      -- CP-element group 279: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1858_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1858_Update/req
      -- 
    ack_4011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1858_inst_ack_0, ack => convolution3D_CP_1767_elements(279)); -- 
    req_4015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(279), ack => WPIPE_maxpool_output_pipe_1858_inst_req_1); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1858_update_completed_
      -- CP-element group 280: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1858_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1858_Update/ack
      -- 
    ack_4016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1858_inst_ack_1, ack => convolution3D_CP_1767_elements(280)); -- 
    -- CP-element group 281:  join  transition  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	271 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1861_sample_start_
      -- CP-element group 281: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1861_Sample/$entry
      -- CP-element group 281: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1861_Sample/req
      -- 
    req_4024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(281), ack => WPIPE_maxpool_output_pipe_1861_inst_req_0); -- 
    convolution3D_cp_element_group_281: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_281"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(271) & convolution3D_CP_1767_elements(280);
      gj_convolution3D_cp_element_group_281 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(281), clk => clk, reset => reset); --
    end block;
    -- CP-element group 282:  transition  input  output  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (6) 
      -- CP-element group 282: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1861_sample_completed_
      -- CP-element group 282: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1861_update_start_
      -- CP-element group 282: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1861_Sample/$exit
      -- CP-element group 282: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1861_Sample/ack
      -- CP-element group 282: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1861_Update/$entry
      -- CP-element group 282: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1861_Update/req
      -- 
    ack_4025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1861_inst_ack_0, ack => convolution3D_CP_1767_elements(282)); -- 
    req_4029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(282), ack => WPIPE_maxpool_output_pipe_1861_inst_req_1); -- 
    -- CP-element group 283:  transition  input  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1861_update_completed_
      -- CP-element group 283: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1861_Update/$exit
      -- CP-element group 283: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1861_Update/ack
      -- 
    ack_4030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1861_inst_ack_1, ack => convolution3D_CP_1767_elements(283)); -- 
    -- CP-element group 284:  join  transition  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	269 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1864_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1864_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1864_Sample/req
      -- 
    req_4038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(284), ack => WPIPE_maxpool_output_pipe_1864_inst_req_0); -- 
    convolution3D_cp_element_group_284: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_284"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(269) & convolution3D_CP_1767_elements(283);
      gj_convolution3D_cp_element_group_284 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(284), clk => clk, reset => reset); --
    end block;
    -- CP-element group 285:  transition  input  output  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	286 
    -- CP-element group 285:  members (6) 
      -- CP-element group 285: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1864_sample_completed_
      -- CP-element group 285: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1864_update_start_
      -- CP-element group 285: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1864_Sample/$exit
      -- CP-element group 285: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1864_Sample/ack
      -- CP-element group 285: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1864_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1864_Update/req
      -- 
    ack_4039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1864_inst_ack_0, ack => convolution3D_CP_1767_elements(285)); -- 
    req_4043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(285), ack => WPIPE_maxpool_output_pipe_1864_inst_req_1); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	285 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1864_update_completed_
      -- CP-element group 286: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1864_Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1864_Update/ack
      -- 
    ack_4044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1864_inst_ack_1, ack => convolution3D_CP_1767_elements(286)); -- 
    -- CP-element group 287:  join  transition  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	267 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1867_sample_start_
      -- CP-element group 287: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1867_Sample/$entry
      -- CP-element group 287: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1867_Sample/req
      -- 
    req_4052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(287), ack => WPIPE_maxpool_output_pipe_1867_inst_req_0); -- 
    convolution3D_cp_element_group_287: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_287"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(267) & convolution3D_CP_1767_elements(286);
      gj_convolution3D_cp_element_group_287 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(287), clk => clk, reset => reset); --
    end block;
    -- CP-element group 288:  transition  input  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (6) 
      -- CP-element group 288: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1867_sample_completed_
      -- CP-element group 288: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1867_update_start_
      -- CP-element group 288: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1867_Sample/$exit
      -- CP-element group 288: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1867_Sample/ack
      -- CP-element group 288: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1867_Update/$entry
      -- CP-element group 288: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1867_Update/req
      -- 
    ack_4053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1867_inst_ack_0, ack => convolution3D_CP_1767_elements(288)); -- 
    req_4057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(288), ack => WPIPE_maxpool_output_pipe_1867_inst_req_1); -- 
    -- CP-element group 289:  transition  input  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1867_update_completed_
      -- CP-element group 289: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1867_Update/$exit
      -- CP-element group 289: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1867_Update/ack
      -- 
    ack_4058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1867_inst_ack_1, ack => convolution3D_CP_1767_elements(289)); -- 
    -- CP-element group 290:  join  transition  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	265 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1870_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1870_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1870_Sample/req
      -- 
    req_4066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(290), ack => WPIPE_maxpool_output_pipe_1870_inst_req_0); -- 
    convolution3D_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(265) & convolution3D_CP_1767_elements(289);
      gj_convolution3D_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1870_sample_completed_
      -- CP-element group 291: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1870_update_start_
      -- CP-element group 291: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1870_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1870_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1870_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1870_Update/req
      -- 
    ack_4067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1870_inst_ack_0, ack => convolution3D_CP_1767_elements(291)); -- 
    req_4071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(291), ack => WPIPE_maxpool_output_pipe_1870_inst_req_1); -- 
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1870_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1870_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1870_Update/ack
      -- 
    ack_4072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1870_inst_ack_1, ack => convolution3D_CP_1767_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: 	263 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1873_sample_start_
      -- CP-element group 293: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1873_Sample/$entry
      -- CP-element group 293: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1873_Sample/req
      -- 
    req_4080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(293), ack => WPIPE_maxpool_output_pipe_1873_inst_req_0); -- 
    convolution3D_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(292) & convolution3D_CP_1767_elements(263);
      gj_convolution3D_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1873_sample_completed_
      -- CP-element group 294: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1873_update_start_
      -- CP-element group 294: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1873_Sample/$exit
      -- CP-element group 294: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1873_Sample/ack
      -- CP-element group 294: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1873_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1873_Update/req
      -- 
    ack_4081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1873_inst_ack_0, ack => convolution3D_CP_1767_elements(294)); -- 
    req_4085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(294), ack => WPIPE_maxpool_output_pipe_1873_inst_req_1); -- 
    -- CP-element group 295:  transition  input  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1873_update_completed_
      -- CP-element group 295: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1873_Update/$exit
      -- CP-element group 295: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1873_Update/ack
      -- 
    ack_4086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1873_inst_ack_1, ack => convolution3D_CP_1767_elements(295)); -- 
    -- CP-element group 296:  join  transition  output  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: 	261 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1876_sample_start_
      -- CP-element group 296: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1876_Sample/$entry
      -- CP-element group 296: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1876_Sample/req
      -- 
    req_4094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(296), ack => WPIPE_maxpool_output_pipe_1876_inst_req_0); -- 
    convolution3D_cp_element_group_296: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_296"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(295) & convolution3D_CP_1767_elements(261);
      gj_convolution3D_cp_element_group_296 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(296), clk => clk, reset => reset); --
    end block;
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1876_sample_completed_
      -- CP-element group 297: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1876_update_start_
      -- CP-element group 297: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1876_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1876_Sample/ack
      -- CP-element group 297: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1876_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1876_Update/req
      -- 
    ack_4095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1876_inst_ack_0, ack => convolution3D_CP_1767_elements(297)); -- 
    req_4099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(297), ack => WPIPE_maxpool_output_pipe_1876_inst_req_1); -- 
    -- CP-element group 298:  transition  place  input  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298:  members (16) 
      -- CP-element group 298: 	 branch_block_stmt_554/branch_block_stmt_554__exit__
      -- CP-element group 298: 	 branch_block_stmt_554/$exit
      -- CP-element group 298: 	 $exit
      -- CP-element group 298: 	 branch_block_stmt_554/merge_stmt_1881__exit__
      -- CP-element group 298: 	 branch_block_stmt_554/return__
      -- CP-element group 298: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878__exit__
      -- CP-element group 298: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/$exit
      -- CP-element group 298: 	 branch_block_stmt_554/merge_stmt_1881_PhiReqMerge
      -- CP-element group 298: 	 branch_block_stmt_554/return___PhiReq/$entry
      -- CP-element group 298: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1876_update_completed_
      -- CP-element group 298: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1876_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_554/call_stmt_1770_to_assign_stmt_1878/WPIPE_maxpool_output_pipe_1876_Update/ack
      -- CP-element group 298: 	 branch_block_stmt_554/merge_stmt_1881_PhiAck/dummy
      -- CP-element group 298: 	 branch_block_stmt_554/merge_stmt_1881_PhiAck/$exit
      -- CP-element group 298: 	 branch_block_stmt_554/merge_stmt_1881_PhiAck/$entry
      -- CP-element group 298: 	 branch_block_stmt_554/return___PhiReq/$exit
      -- 
    ack_4100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1876_inst_ack_1, ack => convolution3D_CP_1767_elements(298)); -- 
    -- CP-element group 299:  transition  output  delay-element  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	86 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	303 
    -- CP-element group 299:  members (5) 
      -- CP-element group 299: 	 branch_block_stmt_554/bbx_xnph369_forx_xbody_PhiReq/$exit
      -- CP-element group 299: 	 branch_block_stmt_554/bbx_xnph369_forx_xbody_PhiReq/phi_stmt_864/$exit
      -- CP-element group 299: 	 branch_block_stmt_554/bbx_xnph369_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_sources/$exit
      -- CP-element group 299: 	 branch_block_stmt_554/bbx_xnph369_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_sources/type_cast_868_konst_delay_trans
      -- CP-element group 299: 	 branch_block_stmt_554/bbx_xnph369_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_req
      -- 
    phi_stmt_864_req_4123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_864_req_4123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(299), ack => phi_stmt_864_req_0); -- 
    -- Element group convolution3D_CP_1767_elements(299) is a control-delay.
    cp_element_299_delay: control_delay_element  generic map(name => " 299_delay", delay_value => 1)  port map(req => convolution3D_CP_1767_elements(86), ack => convolution3D_CP_1767_elements(299), clk => clk, reset =>reset);
    -- CP-element group 300:  transition  input  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	128 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	302 
    -- CP-element group 300:  members (2) 
      -- CP-element group 300: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_sources/type_cast_870/SplitProtocol/Sample/$exit
      -- CP-element group 300: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_sources/type_cast_870/SplitProtocol/Sample/ra
      -- 
    ra_4143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_870_inst_ack_0, ack => convolution3D_CP_1767_elements(300)); -- 
    -- CP-element group 301:  transition  input  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	128 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (2) 
      -- CP-element group 301: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_sources/type_cast_870/SplitProtocol/Update/$exit
      -- CP-element group 301: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_sources/type_cast_870/SplitProtocol/Update/ca
      -- 
    ca_4148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_870_inst_ack_1, ack => convolution3D_CP_1767_elements(301)); -- 
    -- CP-element group 302:  join  transition  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	300 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (6) 
      -- CP-element group 302: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 302: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/phi_stmt_864/$exit
      -- CP-element group 302: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_sources/$exit
      -- CP-element group 302: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_sources/type_cast_870/$exit
      -- CP-element group 302: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_sources/type_cast_870/SplitProtocol/$exit
      -- CP-element group 302: 	 branch_block_stmt_554/forx_xbody_forx_xbody_PhiReq/phi_stmt_864/phi_stmt_864_req
      -- 
    phi_stmt_864_req_4149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_864_req_4149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(302), ack => phi_stmt_864_req_1); -- 
    convolution3D_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(300) & convolution3D_CP_1767_elements(301);
      gj_convolution3D_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  merge  transition  place  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	299 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (2) 
      -- CP-element group 303: 	 branch_block_stmt_554/merge_stmt_863_PhiReqMerge
      -- CP-element group 303: 	 branch_block_stmt_554/merge_stmt_863_PhiAck/$entry
      -- 
    convolution3D_CP_1767_elements(303) <= OrReduce(convolution3D_CP_1767_elements(299) & convolution3D_CP_1767_elements(302));
    -- CP-element group 304:  fork  transition  place  input  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	106 
    -- CP-element group 304: 	110 
    -- CP-element group 304: 	118 
    -- CP-element group 304: 	122 
    -- CP-element group 304: 	114 
    -- CP-element group 304: 	125 
    -- CP-element group 304: 	87 
    -- CP-element group 304: 	88 
    -- CP-element group 304: 	90 
    -- CP-element group 304: 	91 
    -- CP-element group 304: 	94 
    -- CP-element group 304: 	98 
    -- CP-element group 304: 	102 
    -- CP-element group 304:  members (56) 
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_884_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_index_scale_1/scale_rename_ack
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_final_index_sum_regn_Sample/req
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_index_computed_1
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_884_Update/cr
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_933_update_start_
      -- CP-element group 304: 	 branch_block_stmt_554/merge_stmt_863__exit__
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_index_resize_1/index_resize_ack
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026__entry__
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_final_index_sum_regn_update_start
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_1005_update_start_
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_index_scaled_1
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/addr_of_877_complete/$entry
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_969_update_start_
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_index_scale_1/scale_rename_req
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_final_index_sum_regn_Update/req
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_969_Update/cr
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_final_index_sum_regn_Sample/$entry
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Update/word_access_complete/$entry
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_index_resize_1/$entry
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_933_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_index_resize_1/index_resize_req
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_index_resize_1/$exit
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_index_scale_1/$entry
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_index_scale_1/$exit
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_915_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_969_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_915_Update/cr
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_final_index_sum_regn_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Update/word_access_complete/word_0/cr
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_884_update_start_
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_915_update_start_
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_987_Update/cr
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_987_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_Update/word_access_complete/word_0/$entry
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_951_Update/cr
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_951_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_987_update_start_
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_951_update_start_
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/array_obj_ref_876_index_resized_1
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/ptr_deref_1013_update_start_
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_897_Update/cr
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_880_Sample/rr
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_1005_Update/cr
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_880_Sample/$entry
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_897_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_1005_Update/$entry
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_897_update_start_
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/RPIPE_maxpool_input_pipe_880_sample_start_
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/addr_of_877_complete/req
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/type_cast_933_Update/cr
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/$entry
      -- CP-element group 304: 	 branch_block_stmt_554/assign_stmt_878_to_assign_stmt_1026/addr_of_877_update_start_
      -- CP-element group 304: 	 branch_block_stmt_554/merge_stmt_863_PhiAck/$exit
      -- CP-element group 304: 	 branch_block_stmt_554/merge_stmt_863_PhiAck/phi_stmt_864_ack
      -- 
    phi_stmt_864_ack_4154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_864_ack_0, ack => convolution3D_CP_1767_elements(304)); -- 
    req_2471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(304), ack => array_obj_ref_876_index_offset_req_0); -- 
    cr_2519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(304), ack => type_cast_884_inst_req_1); -- 
    req_2476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(304), ack => array_obj_ref_876_index_offset_req_1); -- 
    cr_2659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(304), ack => type_cast_969_inst_req_1); -- 
    cr_2575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(304), ack => type_cast_915_inst_req_1); -- 
    cr_2765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(304), ack => ptr_deref_1013_store_0_req_1); -- 
    cr_2687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(304), ack => type_cast_987_inst_req_1); -- 
    cr_2631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(304), ack => type_cast_951_inst_req_1); -- 
    cr_2547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(304), ack => type_cast_897_inst_req_1); -- 
    rr_2500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(304), ack => RPIPE_maxpool_input_pipe_880_inst_req_0); -- 
    cr_2715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(304), ack => type_cast_1005_inst_req_1); -- 
    req_2491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(304), ack => addr_of_877_final_reg_req_1); -- 
    cr_2603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(304), ack => type_cast_933_inst_req_1); -- 
    -- CP-element group 305:  transition  output  delay-element  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	76 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	309 
    -- CP-element group 305:  members (5) 
      -- CP-element group 305: 	 branch_block_stmt_554/entry_forx_xend_PhiReq/$exit
      -- CP-element group 305: 	 branch_block_stmt_554/entry_forx_xend_PhiReq/phi_stmt_1058/$exit
      -- CP-element group 305: 	 branch_block_stmt_554/entry_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_sources/$exit
      -- CP-element group 305: 	 branch_block_stmt_554/entry_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_sources/type_cast_1064_konst_delay_trans
      -- CP-element group 305: 	 branch_block_stmt_554/entry_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_req
      -- 
    phi_stmt_1058_req_4177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1058_req_4177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(305), ack => phi_stmt_1058_req_1); -- 
    -- Element group convolution3D_CP_1767_elements(305) is a control-delay.
    cp_element_305_delay: control_delay_element  generic map(name => " 305_delay", delay_value => 1)  port map(req => convolution3D_CP_1767_elements(76), ack => convolution3D_CP_1767_elements(305), clk => clk, reset =>reset);
    -- CP-element group 306:  transition  input  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	127 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	308 
    -- CP-element group 306:  members (2) 
      -- CP-element group 306: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_sources/type_cast_1061/SplitProtocol/Sample/$exit
      -- CP-element group 306: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_sources/type_cast_1061/SplitProtocol/Sample/ra
      -- 
    ra_4197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1061_inst_ack_0, ack => convolution3D_CP_1767_elements(306)); -- 
    -- CP-element group 307:  transition  input  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	127 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (2) 
      -- CP-element group 307: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_sources/type_cast_1061/SplitProtocol/Update/$exit
      -- CP-element group 307: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_sources/type_cast_1061/SplitProtocol/Update/ca
      -- 
    ca_4202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1061_inst_ack_1, ack => convolution3D_CP_1767_elements(307)); -- 
    -- CP-element group 308:  join  transition  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	306 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (6) 
      -- CP-element group 308: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$exit
      -- CP-element group 308: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1058/$exit
      -- CP-element group 308: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_sources/$exit
      -- CP-element group 308: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_sources/type_cast_1061/$exit
      -- CP-element group 308: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_sources/type_cast_1061/SplitProtocol/$exit
      -- CP-element group 308: 	 branch_block_stmt_554/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1058/phi_stmt_1058_req
      -- 
    phi_stmt_1058_req_4203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1058_req_4203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(308), ack => phi_stmt_1058_req_0); -- 
    convolution3D_cp_element_group_308: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_308"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(306) & convolution3D_CP_1767_elements(307);
      gj_convolution3D_cp_element_group_308 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(308), clk => clk, reset => reset); --
    end block;
    -- CP-element group 309:  merge  transition  place  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	305 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (2) 
      -- CP-element group 309: 	 branch_block_stmt_554/merge_stmt_1057_PhiReqMerge
      -- CP-element group 309: 	 branch_block_stmt_554/merge_stmt_1057_PhiAck/$entry
      -- 
    convolution3D_CP_1767_elements(309) <= OrReduce(convolution3D_CP_1767_elements(305) & convolution3D_CP_1767_elements(308));
    -- CP-element group 310:  branch  transition  place  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	129 
    -- CP-element group 310: 	130 
    -- CP-element group 310:  members (15) 
      -- CP-element group 310: 	 branch_block_stmt_554/merge_stmt_1057__exit__
      -- CP-element group 310: 	 branch_block_stmt_554/if_stmt_1078_else_link/$entry
      -- CP-element group 310: 	 branch_block_stmt_554/assign_stmt_1071_to_assign_stmt_1077__exit__
      -- CP-element group 310: 	 branch_block_stmt_554/if_stmt_1078__entry__
      -- CP-element group 310: 	 branch_block_stmt_554/assign_stmt_1071_to_assign_stmt_1077__entry__
      -- CP-element group 310: 	 branch_block_stmt_554/R_tobool_1079_place
      -- CP-element group 310: 	 branch_block_stmt_554/if_stmt_1078_if_link/$entry
      -- CP-element group 310: 	 branch_block_stmt_554/if_stmt_1078_eval_test/branch_req
      -- CP-element group 310: 	 branch_block_stmt_554/if_stmt_1078_eval_test/$exit
      -- CP-element group 310: 	 branch_block_stmt_554/if_stmt_1078_eval_test/$entry
      -- CP-element group 310: 	 branch_block_stmt_554/if_stmt_1078_dead_link/$entry
      -- CP-element group 310: 	 branch_block_stmt_554/assign_stmt_1071_to_assign_stmt_1077/$exit
      -- CP-element group 310: 	 branch_block_stmt_554/assign_stmt_1071_to_assign_stmt_1077/$entry
      -- CP-element group 310: 	 branch_block_stmt_554/merge_stmt_1057_PhiAck/$exit
      -- CP-element group 310: 	 branch_block_stmt_554/merge_stmt_1057_PhiAck/phi_stmt_1058_ack
      -- 
    phi_stmt_1058_ack_4208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1058_ack_0, ack => convolution3D_CP_1767_elements(310)); -- 
    branch_req_2799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(310), ack => if_stmt_1078_branch_req_0); -- 
    -- CP-element group 311:  transition  output  delay-element  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	130 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	313 
    -- CP-element group 311:  members (4) 
      -- CP-element group 311: 	 branch_block_stmt_554/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/$exit
      -- CP-element group 311: 	 branch_block_stmt_554/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_sources/$exit
      -- CP-element group 311: 	 branch_block_stmt_554/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_sources/type_cast_1103_konst_delay_trans
      -- CP-element group 311: 	 branch_block_stmt_554/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_req
      -- 
    phi_stmt_1099_req_4231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1099_req_4231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(311), ack => phi_stmt_1099_req_0); -- 
    -- Element group convolution3D_CP_1767_elements(311) is a control-delay.
    cp_element_311_delay: control_delay_element  generic map(name => " 311_delay", delay_value => 1)  port map(req => convolution3D_CP_1767_elements(130), ack => convolution3D_CP_1767_elements(311), clk => clk, reset =>reset);
    -- CP-element group 312:  transition  output  delay-element  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	130 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (4) 
      -- CP-element group 312: 	 branch_block_stmt_554/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/$exit
      -- CP-element group 312: 	 branch_block_stmt_554/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/$exit
      -- CP-element group 312: 	 branch_block_stmt_554/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1110_konst_delay_trans
      -- CP-element group 312: 	 branch_block_stmt_554/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_req
      -- 
    phi_stmt_1106_req_4239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1106_req_4239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(312), ack => phi_stmt_1106_req_0); -- 
    -- Element group convolution3D_CP_1767_elements(312) is a control-delay.
    cp_element_312_delay: control_delay_element  generic map(name => " 312_delay", delay_value => 1)  port map(req => convolution3D_CP_1767_elements(130), ack => convolution3D_CP_1767_elements(312), clk => clk, reset =>reset);
    -- CP-element group 313:  join  transition  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	311 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	321 
    -- CP-element group 313:  members (1) 
      -- CP-element group 313: 	 branch_block_stmt_554/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_313: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_313"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(311) & convolution3D_CP_1767_elements(312);
      gj_convolution3D_cp_element_group_313 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(313), clk => clk, reset => reset); --
    end block;
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	138 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	316 
    -- CP-element group 314:  members (2) 
      -- CP-element group 314: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_sources/type_cast_1105/SplitProtocol/Sample/$exit
      -- CP-element group 314: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_sources/type_cast_1105/SplitProtocol/Sample/ra
      -- 
    ra_4259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1105_inst_ack_0, ack => convolution3D_CP_1767_elements(314)); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	138 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	316 
    -- CP-element group 315:  members (2) 
      -- CP-element group 315: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_sources/type_cast_1105/SplitProtocol/Update/$exit
      -- CP-element group 315: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_sources/type_cast_1105/SplitProtocol/Update/ca
      -- 
    ca_4264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1105_inst_ack_1, ack => convolution3D_CP_1767_elements(315)); -- 
    -- CP-element group 316:  join  transition  output  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	314 
    -- CP-element group 316: 	315 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	320 
    -- CP-element group 316:  members (5) 
      -- CP-element group 316: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/$exit
      -- CP-element group 316: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_sources/$exit
      -- CP-element group 316: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_sources/type_cast_1105/$exit
      -- CP-element group 316: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_sources/type_cast_1105/SplitProtocol/$exit
      -- CP-element group 316: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1099/phi_stmt_1099_req
      -- 
    phi_stmt_1099_req_4265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1099_req_4265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(316), ack => phi_stmt_1099_req_1); -- 
    convolution3D_cp_element_group_316: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_316"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(314) & convolution3D_CP_1767_elements(315);
      gj_convolution3D_cp_element_group_316 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(316), clk => clk, reset => reset); --
    end block;
    -- CP-element group 317:  transition  input  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	138 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	319 
    -- CP-element group 317:  members (2) 
      -- CP-element group 317: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/Sample/$exit
      -- CP-element group 317: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/Sample/ra
      -- 
    ra_4282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1112_inst_ack_0, ack => convolution3D_CP_1767_elements(317)); -- 
    -- CP-element group 318:  transition  input  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	138 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (2) 
      -- CP-element group 318: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/Update/$exit
      -- CP-element group 318: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/Update/ca
      -- 
    ca_4287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1112_inst_ack_1, ack => convolution3D_CP_1767_elements(318)); -- 
    -- CP-element group 319:  join  transition  output  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	317 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	320 
    -- CP-element group 319:  members (5) 
      -- CP-element group 319: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/$exit
      -- CP-element group 319: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/$exit
      -- CP-element group 319: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/$exit
      -- CP-element group 319: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/$exit
      -- CP-element group 319: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1106/phi_stmt_1106_req
      -- 
    phi_stmt_1106_req_4288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1106_req_4288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(319), ack => phi_stmt_1106_req_1); -- 
    convolution3D_cp_element_group_319: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_319"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(317) & convolution3D_CP_1767_elements(318);
      gj_convolution3D_cp_element_group_319 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(319), clk => clk, reset => reset); --
    end block;
    -- CP-element group 320:  join  transition  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	316 
    -- CP-element group 320: 	319 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	321 
    -- CP-element group 320:  members (1) 
      -- CP-element group 320: 	 branch_block_stmt_554/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_320: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_320"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(316) & convolution3D_CP_1767_elements(319);
      gj_convolution3D_cp_element_group_320 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(320), clk => clk, reset => reset); --
    end block;
    -- CP-element group 321:  merge  fork  transition  place  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	313 
    -- CP-element group 321: 	320 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321: 	323 
    -- CP-element group 321:  members (2) 
      -- CP-element group 321: 	 branch_block_stmt_554/merge_stmt_1098_PhiReqMerge
      -- CP-element group 321: 	 branch_block_stmt_554/merge_stmt_1098_PhiAck/$entry
      -- 
    convolution3D_CP_1767_elements(321) <= OrReduce(convolution3D_CP_1767_elements(313) & convolution3D_CP_1767_elements(320));
    -- CP-element group 322:  transition  input  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	324 
    -- CP-element group 322:  members (1) 
      -- CP-element group 322: 	 branch_block_stmt_554/merge_stmt_1098_PhiAck/phi_stmt_1099_ack
      -- 
    phi_stmt_1099_ack_4293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1099_ack_0, ack => convolution3D_CP_1767_elements(322)); -- 
    -- CP-element group 323:  transition  input  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	321 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (1) 
      -- CP-element group 323: 	 branch_block_stmt_554/merge_stmt_1098_PhiAck/phi_stmt_1106_ack
      -- 
    phi_stmt_1106_ack_4294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1106_ack_0, ack => convolution3D_CP_1767_elements(323)); -- 
    -- CP-element group 324:  join  fork  transition  place  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	322 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	131 
    -- CP-element group 324: 	134 
    -- CP-element group 324: 	135 
    -- CP-element group 324: 	136 
    -- CP-element group 324:  members (16) 
      -- CP-element group 324: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1146_update_start_
      -- CP-element group 324: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152__entry__
      -- CP-element group 324: 	 branch_block_stmt_554/merge_stmt_1098__exit__
      -- CP-element group 324: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1131_Update/$entry
      -- CP-element group 324: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1146_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1131_Update/cr
      -- CP-element group 324: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1131_update_start_
      -- CP-element group 324: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1146_Update/cr
      -- CP-element group 324: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1146_Update/$entry
      -- CP-element group 324: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1146_Sample/rr
      -- CP-element group 324: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/type_cast_1146_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/RPIPE_maxpool_input_pipe_1127_Sample/rr
      -- CP-element group 324: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/RPIPE_maxpool_input_pipe_1127_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/RPIPE_maxpool_input_pipe_1127_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_554/assign_stmt_1119_to_assign_stmt_1152/$entry
      -- CP-element group 324: 	 branch_block_stmt_554/merge_stmt_1098_PhiAck/$exit
      -- 
    cr_2843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(324), ack => type_cast_1131_inst_req_1); -- 
    cr_2857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(324), ack => type_cast_1146_inst_req_1); -- 
    rr_2852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(324), ack => type_cast_1146_inst_req_0); -- 
    rr_2824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(324), ack => RPIPE_maxpool_input_pipe_1127_inst_req_0); -- 
    convolution3D_cp_element_group_324: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_324"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(322) & convolution3D_CP_1767_elements(323);
      gj_convolution3D_cp_element_group_324 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(324), clk => clk, reset => reset); --
    end block;
    -- CP-element group 325:  transition  input  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	139 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	327 
    -- CP-element group 325:  members (2) 
      -- CP-element group 325: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1160/phi_stmt_1160_sources/type_cast_1163/SplitProtocol/Sample/$exit
      -- CP-element group 325: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1160/phi_stmt_1160_sources/type_cast_1163/SplitProtocol/Sample/ra
      -- 
    ra_4318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1163_inst_ack_0, ack => convolution3D_CP_1767_elements(325)); -- 
    -- CP-element group 326:  transition  input  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	139 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (2) 
      -- CP-element group 326: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1160/phi_stmt_1160_sources/type_cast_1163/SplitProtocol/Update/$exit
      -- CP-element group 326: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1160/phi_stmt_1160_sources/type_cast_1163/SplitProtocol/Update/ca
      -- 
    ca_4323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1163_inst_ack_1, ack => convolution3D_CP_1767_elements(326)); -- 
    -- CP-element group 327:  join  transition  place  output  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	325 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327:  members (8) 
      -- CP-element group 327: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$exit
      -- CP-element group 327: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1160/$exit
      -- CP-element group 327: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1160/phi_stmt_1160_sources/$exit
      -- CP-element group 327: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1160/phi_stmt_1160_sources/type_cast_1163/$exit
      -- CP-element group 327: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1160/phi_stmt_1160_sources/type_cast_1163/SplitProtocol/$exit
      -- CP-element group 327: 	 branch_block_stmt_554/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1160/phi_stmt_1160_req
      -- CP-element group 327: 	 branch_block_stmt_554/merge_stmt_1159_PhiReqMerge
      -- CP-element group 327: 	 branch_block_stmt_554/merge_stmt_1159_PhiAck/$entry
      -- 
    phi_stmt_1160_req_4324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1160_req_4324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(327), ack => phi_stmt_1160_req_0); -- 
    convolution3D_cp_element_group_327: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_327"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(325) & convolution3D_CP_1767_elements(326);
      gj_convolution3D_cp_element_group_327 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(327), clk => clk, reset => reset); --
    end block;
    -- CP-element group 328:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	145 
    -- CP-element group 328: 	140 
    -- CP-element group 328: 	141 
    -- CP-element group 328: 	143 
    -- CP-element group 328:  members (29) 
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_index_scale_1/$entry
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_index_computed_1
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_final_index_sum_regn_Sample/req
      -- CP-element group 328: 	 branch_block_stmt_554/merge_stmt_1159__exit__
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198__entry__
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_index_scale_1/scale_rename_ack
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_index_scale_1/scale_rename_req
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_index_resized_1
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_index_scaled_1
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_index_scale_1/$exit
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_index_resize_1/index_resize_ack
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/addr_of_1193_update_start_
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_final_index_sum_regn_update_start
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_final_index_sum_regn_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_index_resize_1/index_resize_req
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_index_resize_1/$entry
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_index_resize_1/$exit
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/$entry
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_final_index_sum_regn_Update/$entry
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/array_obj_ref_1192_final_index_sum_regn_Update/req
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/addr_of_1193_complete/$entry
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/addr_of_1193_complete/req
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_update_start_
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Update/$entry
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Update/word_access_complete/$entry
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Update/word_access_complete/word_0/$entry
      -- CP-element group 328: 	 branch_block_stmt_554/assign_stmt_1170_to_assign_stmt_1198/ptr_deref_1196_Update/word_access_complete/word_0/cr
      -- CP-element group 328: 	 branch_block_stmt_554/merge_stmt_1159_PhiAck/$exit
      -- CP-element group 328: 	 branch_block_stmt_554/merge_stmt_1159_PhiAck/phi_stmt_1160_ack
      -- 
    phi_stmt_1160_ack_4329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1160_ack_0, ack => convolution3D_CP_1767_elements(328)); -- 
    req_2905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(328), ack => array_obj_ref_1192_index_offset_req_0); -- 
    req_2910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(328), ack => array_obj_ref_1192_index_offset_req_1); -- 
    req_2925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(328), ack => addr_of_1193_final_reg_req_1); -- 
    cr_2975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(328), ack => ptr_deref_1196_store_0_req_1); -- 
    -- CP-element group 329:  merge  fork  transition  place  output  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	146 
    -- CP-element group 329: 	129 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	147 
    -- CP-element group 329: 	148 
    -- CP-element group 329: 	149 
    -- CP-element group 329: 	150 
    -- CP-element group 329: 	151 
    -- CP-element group 329: 	152 
    -- CP-element group 329:  members (25) 
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248__entry__
      -- CP-element group 329: 	 branch_block_stmt_554/merge_stmt_1200__exit__
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/$entry
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1203_sample_start_
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1203_update_start_
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1203_Sample/$entry
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1203_Sample/rr
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1203_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1203_Update/cr
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1207_sample_start_
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1207_update_start_
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1207_Sample/$entry
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1207_Sample/rr
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1207_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1207_Update/cr
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1211_sample_start_
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1211_update_start_
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1211_Sample/$entry
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1211_Sample/rr
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1211_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_554/assign_stmt_1204_to_assign_stmt_1248/type_cast_1211_Update/cr
      -- CP-element group 329: 	 branch_block_stmt_554/merge_stmt_1200_PhiReqMerge
      -- CP-element group 329: 	 branch_block_stmt_554/merge_stmt_1200_PhiAck/$entry
      -- CP-element group 329: 	 branch_block_stmt_554/merge_stmt_1200_PhiAck/$exit
      -- CP-element group 329: 	 branch_block_stmt_554/merge_stmt_1200_PhiAck/dummy
      -- 
    rr_2987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(329), ack => type_cast_1203_inst_req_0); -- 
    cr_2992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(329), ack => type_cast_1203_inst_req_1); -- 
    rr_3001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(329), ack => type_cast_1207_inst_req_0); -- 
    cr_3006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(329), ack => type_cast_1207_inst_req_1); -- 
    rr_3015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(329), ack => type_cast_1211_inst_req_0); -- 
    cr_3020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(329), ack => type_cast_1211_inst_req_1); -- 
    convolution3D_CP_1767_elements(329) <= OrReduce(convolution3D_CP_1767_elements(146) & convolution3D_CP_1767_elements(129));
    -- CP-element group 330:  transition  output  delay-element  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	166 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	334 
    -- CP-element group 330:  members (5) 
      -- CP-element group 330: 	 branch_block_stmt_554/bbx_xnph_forx_xbody163_PhiReq/$exit
      -- CP-element group 330: 	 branch_block_stmt_554/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1325/$exit
      -- CP-element group 330: 	 branch_block_stmt_554/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_sources/$exit
      -- CP-element group 330: 	 branch_block_stmt_554/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_sources/type_cast_1329_konst_delay_trans
      -- CP-element group 330: 	 branch_block_stmt_554/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_req
      -- 
    phi_stmt_1325_req_4363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1325_req_4363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(330), ack => phi_stmt_1325_req_0); -- 
    -- Element group convolution3D_CP_1767_elements(330) is a control-delay.
    cp_element_330_delay: control_delay_element  generic map(name => " 330_delay", delay_value => 1)  port map(req => convolution3D_CP_1767_elements(166), ack => convolution3D_CP_1767_elements(330), clk => clk, reset =>reset);
    -- CP-element group 331:  transition  input  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	208 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	333 
    -- CP-element group 331:  members (2) 
      -- CP-element group 331: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_sources/type_cast_1331/SplitProtocol/Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_sources/type_cast_1331/SplitProtocol/Sample/ra
      -- 
    ra_4383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1331_inst_ack_0, ack => convolution3D_CP_1767_elements(331)); -- 
    -- CP-element group 332:  transition  input  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	208 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (2) 
      -- CP-element group 332: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_sources/type_cast_1331/SplitProtocol/Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_sources/type_cast_1331/SplitProtocol/Update/ca
      -- 
    ca_4388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1331_inst_ack_1, ack => convolution3D_CP_1767_elements(332)); -- 
    -- CP-element group 333:  join  transition  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	331 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (6) 
      -- CP-element group 333: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/$exit
      -- CP-element group 333: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1325/$exit
      -- CP-element group 333: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_sources/$exit
      -- CP-element group 333: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_sources/type_cast_1331/$exit
      -- CP-element group 333: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_sources/type_cast_1331/SplitProtocol/$exit
      -- CP-element group 333: 	 branch_block_stmt_554/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1325/phi_stmt_1325_req
      -- 
    phi_stmt_1325_req_4389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1325_req_4389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(333), ack => phi_stmt_1325_req_1); -- 
    convolution3D_cp_element_group_333: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_333"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(331) & convolution3D_CP_1767_elements(332);
      gj_convolution3D_cp_element_group_333 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(333), clk => clk, reset => reset); --
    end block;
    -- CP-element group 334:  merge  transition  place  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	330 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (2) 
      -- CP-element group 334: 	 branch_block_stmt_554/merge_stmt_1324_PhiReqMerge
      -- CP-element group 334: 	 branch_block_stmt_554/merge_stmt_1324_PhiAck/$entry
      -- 
    convolution3D_CP_1767_elements(334) <= OrReduce(convolution3D_CP_1767_elements(330) & convolution3D_CP_1767_elements(333));
    -- CP-element group 335:  fork  transition  place  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	167 
    -- CP-element group 335: 	186 
    -- CP-element group 335: 	168 
    -- CP-element group 335: 	170 
    -- CP-element group 335: 	182 
    -- CP-element group 335: 	205 
    -- CP-element group 335: 	171 
    -- CP-element group 335: 	174 
    -- CP-element group 335: 	178 
    -- CP-element group 335: 	190 
    -- CP-element group 335: 	194 
    -- CP-element group 335: 	198 
    -- CP-element group 335: 	202 
    -- CP-element group 335:  members (56) 
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487__entry__
      -- CP-element group 335: 	 branch_block_stmt_554/merge_stmt_1324__exit__
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/$entry
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/addr_of_1338_update_start_
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_index_resized_1
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_index_scaled_1
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_index_computed_1
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_index_resize_1/$entry
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_index_resize_1/$exit
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_index_resize_1/index_resize_req
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_index_resize_1/index_resize_ack
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_index_scale_1/$entry
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_index_scale_1/$exit
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_index_scale_1/scale_rename_req
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_index_scale_1/scale_rename_ack
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_final_index_sum_regn_update_start
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_final_index_sum_regn_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_final_index_sum_regn_Sample/req
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_final_index_sum_regn_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/array_obj_ref_1337_final_index_sum_regn_Update/req
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/addr_of_1338_complete/$entry
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/addr_of_1338_complete/req
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1341_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1341_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/RPIPE_maxpool_input_pipe_1341_Sample/rr
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1345_update_start_
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1345_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1345_Update/cr
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1358_update_start_
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1358_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1358_Update/cr
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1376_update_start_
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1376_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1376_Update/cr
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1394_update_start_
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1394_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1394_Update/cr
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1412_update_start_
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1412_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1412_Update/cr
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1430_update_start_
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1430_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1430_Update/cr
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1448_update_start_
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1448_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1448_Update/cr
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1466_update_start_
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1466_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/type_cast_1466_Update/cr
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_update_start_
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Update/word_access_complete/$entry
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Update/word_access_complete/word_0/$entry
      -- CP-element group 335: 	 branch_block_stmt_554/assign_stmt_1339_to_assign_stmt_1487/ptr_deref_1474_Update/word_access_complete/word_0/cr
      -- CP-element group 335: 	 branch_block_stmt_554/merge_stmt_1324_PhiAck/$exit
      -- CP-element group 335: 	 branch_block_stmt_554/merge_stmt_1324_PhiAck/phi_stmt_1325_ack
      -- 
    phi_stmt_1325_ack_4394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1325_ack_0, ack => convolution3D_CP_1767_elements(335)); -- 
    req_3141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(335), ack => array_obj_ref_1337_index_offset_req_0); -- 
    req_3146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(335), ack => array_obj_ref_1337_index_offset_req_1); -- 
    req_3161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(335), ack => addr_of_1338_final_reg_req_1); -- 
    rr_3170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(335), ack => RPIPE_maxpool_input_pipe_1341_inst_req_0); -- 
    cr_3189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(335), ack => type_cast_1345_inst_req_1); -- 
    cr_3217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(335), ack => type_cast_1358_inst_req_1); -- 
    cr_3245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(335), ack => type_cast_1376_inst_req_1); -- 
    cr_3273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(335), ack => type_cast_1394_inst_req_1); -- 
    cr_3301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(335), ack => type_cast_1412_inst_req_1); -- 
    cr_3329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(335), ack => type_cast_1430_inst_req_1); -- 
    cr_3357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(335), ack => type_cast_1448_inst_req_1); -- 
    cr_3385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(335), ack => type_cast_1466_inst_req_1); -- 
    cr_3435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(335), ack => ptr_deref_1474_store_0_req_1); -- 
    -- CP-element group 336:  transition  input  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	207 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	338 
    -- CP-element group 336:  members (2) 
      -- CP-element group 336: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/Sample/$exit
      -- CP-element group 336: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/Sample/ra
      -- 
    ra_4426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1522_inst_ack_0, ack => convolution3D_CP_1767_elements(336)); -- 
    -- CP-element group 337:  transition  input  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	207 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (2) 
      -- CP-element group 337: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/Update/$exit
      -- CP-element group 337: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/Update/ca
      -- 
    ca_4431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1522_inst_ack_1, ack => convolution3D_CP_1767_elements(337)); -- 
    -- CP-element group 338:  join  transition  output  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	336 
    -- CP-element group 338: 	337 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	340 
    -- CP-element group 338:  members (6) 
      -- CP-element group 338: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/$exit
      -- CP-element group 338: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1519/$exit
      -- CP-element group 338: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/$exit
      -- CP-element group 338: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/$exit
      -- CP-element group 338: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/$exit
      -- CP-element group 338: 	 branch_block_stmt_554/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_req
      -- 
    phi_stmt_1519_req_4432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1519_req_4432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(338), ack => phi_stmt_1519_req_0); -- 
    convolution3D_cp_element_group_338: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_338"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(336) & convolution3D_CP_1767_elements(337);
      gj_convolution3D_cp_element_group_338 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(338), clk => clk, reset => reset); --
    end block;
    -- CP-element group 339:  transition  output  delay-element  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	155 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (5) 
      -- CP-element group 339: 	 branch_block_stmt_554/ifx_xend_forx_xend215_PhiReq/$exit
      -- CP-element group 339: 	 branch_block_stmt_554/ifx_xend_forx_xend215_PhiReq/phi_stmt_1519/$exit
      -- CP-element group 339: 	 branch_block_stmt_554/ifx_xend_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/$exit
      -- CP-element group 339: 	 branch_block_stmt_554/ifx_xend_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1525_konst_delay_trans
      -- CP-element group 339: 	 branch_block_stmt_554/ifx_xend_forx_xend215_PhiReq/phi_stmt_1519/phi_stmt_1519_req
      -- 
    phi_stmt_1519_req_4443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1519_req_4443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(339), ack => phi_stmt_1519_req_1); -- 
    -- Element group convolution3D_CP_1767_elements(339) is a control-delay.
    cp_element_339_delay: control_delay_element  generic map(name => " 339_delay", delay_value => 1)  port map(req => convolution3D_CP_1767_elements(155), ack => convolution3D_CP_1767_elements(339), clk => clk, reset =>reset);
    -- CP-element group 340:  merge  transition  place  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (2) 
      -- CP-element group 340: 	 branch_block_stmt_554/merge_stmt_1518_PhiReqMerge
      -- CP-element group 340: 	 branch_block_stmt_554/merge_stmt_1518_PhiAck/$entry
      -- 
    convolution3D_CP_1767_elements(340) <= OrReduce(convolution3D_CP_1767_elements(338) & convolution3D_CP_1767_elements(339));
    -- CP-element group 341:  branch  transition  place  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	209 
    -- CP-element group 341: 	210 
    -- CP-element group 341:  members (15) 
      -- CP-element group 341: 	 branch_block_stmt_554/merge_stmt_1518__exit__
      -- CP-element group 341: 	 branch_block_stmt_554/assign_stmt_1532_to_assign_stmt_1538__entry__
      -- CP-element group 341: 	 branch_block_stmt_554/assign_stmt_1532_to_assign_stmt_1538__exit__
      -- CP-element group 341: 	 branch_block_stmt_554/if_stmt_1539__entry__
      -- CP-element group 341: 	 branch_block_stmt_554/assign_stmt_1532_to_assign_stmt_1538/$entry
      -- CP-element group 341: 	 branch_block_stmt_554/assign_stmt_1532_to_assign_stmt_1538/$exit
      -- CP-element group 341: 	 branch_block_stmt_554/if_stmt_1539_dead_link/$entry
      -- CP-element group 341: 	 branch_block_stmt_554/if_stmt_1539_else_link/$entry
      -- CP-element group 341: 	 branch_block_stmt_554/R_tobool218_1540_place
      -- CP-element group 341: 	 branch_block_stmt_554/if_stmt_1539_if_link/$entry
      -- CP-element group 341: 	 branch_block_stmt_554/if_stmt_1539_eval_test/branch_req
      -- CP-element group 341: 	 branch_block_stmt_554/if_stmt_1539_eval_test/$exit
      -- CP-element group 341: 	 branch_block_stmt_554/if_stmt_1539_eval_test/$entry
      -- CP-element group 341: 	 branch_block_stmt_554/merge_stmt_1518_PhiAck/$exit
      -- CP-element group 341: 	 branch_block_stmt_554/merge_stmt_1518_PhiAck/phi_stmt_1519_ack
      -- 
    phi_stmt_1519_ack_4448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1519_ack_0, ack => convolution3D_CP_1767_elements(341)); -- 
    branch_req_3469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(341), ack => if_stmt_1539_branch_req_0); -- 
    -- CP-element group 342:  transition  output  delay-element  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	212 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	344 
    -- CP-element group 342:  members (4) 
      -- CP-element group 342: 	 branch_block_stmt_554/bbx_xnphx_xi340_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/$exit
      -- CP-element group 342: 	 branch_block_stmt_554/bbx_xnphx_xi340_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/$exit
      -- CP-element group 342: 	 branch_block_stmt_554/bbx_xnphx_xi340_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1568_konst_delay_trans
      -- CP-element group 342: 	 branch_block_stmt_554/bbx_xnphx_xi340_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_req
      -- 
    phi_stmt_1564_req_4471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1564_req_4471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(342), ack => phi_stmt_1564_req_0); -- 
    -- Element group convolution3D_CP_1767_elements(342) is a control-delay.
    cp_element_342_delay: control_delay_element  generic map(name => " 342_delay", delay_value => 1)  port map(req => convolution3D_CP_1767_elements(212), ack => convolution3D_CP_1767_elements(342), clk => clk, reset =>reset);
    -- CP-element group 343:  transition  output  delay-element  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	212 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (4) 
      -- CP-element group 343: 	 branch_block_stmt_554/bbx_xnphx_xi340_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_req
      -- CP-element group 343: 	 branch_block_stmt_554/bbx_xnphx_xi340_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_sources/type_cast_1575_konst_delay_trans
      -- CP-element group 343: 	 branch_block_stmt_554/bbx_xnphx_xi340_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/$exit
      -- CP-element group 343: 	 branch_block_stmt_554/bbx_xnphx_xi340_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_sources/$exit
      -- 
    phi_stmt_1571_req_4479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1571_req_4479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(343), ack => phi_stmt_1571_req_0); -- 
    -- Element group convolution3D_CP_1767_elements(343) is a control-delay.
    cp_element_343_delay: control_delay_element  generic map(name => " 343_delay", delay_value => 1)  port map(req => convolution3D_CP_1767_elements(212), ack => convolution3D_CP_1767_elements(343), clk => clk, reset =>reset);
    -- CP-element group 344:  join  transition  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	352 
    -- CP-element group 344:  members (1) 
      -- CP-element group 344: 	 branch_block_stmt_554/bbx_xnphx_xi340_forx_xbodyx_xi349_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_344: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_344"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(342) & convolution3D_CP_1767_elements(343);
      gj_convolution3D_cp_element_group_344 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(344), clk => clk, reset => reset); --
    end block;
    -- CP-element group 345:  transition  input  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	220 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	347 
    -- CP-element group 345:  members (2) 
      -- CP-element group 345: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1570/SplitProtocol/Sample/ra
      -- CP-element group 345: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1570/SplitProtocol/Sample/$exit
      -- 
    ra_4499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1570_inst_ack_0, ack => convolution3D_CP_1767_elements(345)); -- 
    -- CP-element group 346:  transition  input  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	220 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (2) 
      -- CP-element group 346: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1570/SplitProtocol/Update/ca
      -- CP-element group 346: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1570/SplitProtocol/Update/$exit
      -- 
    ca_4504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1570_inst_ack_1, ack => convolution3D_CP_1767_elements(346)); -- 
    -- CP-element group 347:  join  transition  output  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	345 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	351 
    -- CP-element group 347:  members (5) 
      -- CP-element group 347: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1570/SplitProtocol/$exit
      -- CP-element group 347: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/type_cast_1570/$exit
      -- CP-element group 347: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_sources/$exit
      -- CP-element group 347: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/$exit
      -- CP-element group 347: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1564/phi_stmt_1564_req
      -- 
    phi_stmt_1564_req_4505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1564_req_4505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(347), ack => phi_stmt_1564_req_1); -- 
    convolution3D_cp_element_group_347: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_347"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(345) & convolution3D_CP_1767_elements(346);
      gj_convolution3D_cp_element_group_347 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(347), clk => clk, reset => reset); --
    end block;
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	220 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	350 
    -- CP-element group 348:  members (2) 
      -- CP-element group 348: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_sources/type_cast_1577/SplitProtocol/Sample/ra
      -- CP-element group 348: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_sources/type_cast_1577/SplitProtocol/Sample/$exit
      -- 
    ra_4522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1577_inst_ack_0, ack => convolution3D_CP_1767_elements(348)); -- 
    -- CP-element group 349:  transition  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	220 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	350 
    -- CP-element group 349:  members (2) 
      -- CP-element group 349: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_sources/type_cast_1577/SplitProtocol/Update/ca
      -- CP-element group 349: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_sources/type_cast_1577/SplitProtocol/Update/$exit
      -- 
    ca_4527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1577_inst_ack_1, ack => convolution3D_CP_1767_elements(349)); -- 
    -- CP-element group 350:  join  transition  output  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	348 
    -- CP-element group 350: 	349 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	351 
    -- CP-element group 350:  members (5) 
      -- CP-element group 350: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_sources/type_cast_1577/SplitProtocol/$exit
      -- CP-element group 350: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_sources/type_cast_1577/$exit
      -- CP-element group 350: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_sources/$exit
      -- CP-element group 350: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/$exit
      -- CP-element group 350: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/phi_stmt_1571/phi_stmt_1571_req
      -- 
    phi_stmt_1571_req_4528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1571_req_4528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(350), ack => phi_stmt_1571_req_1); -- 
    convolution3D_cp_element_group_350: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_350"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(348) & convolution3D_CP_1767_elements(349);
      gj_convolution3D_cp_element_group_350 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(350), clk => clk, reset => reset); --
    end block;
    -- CP-element group 351:  join  transition  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	347 
    -- CP-element group 351: 	350 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (1) 
      -- CP-element group 351: 	 branch_block_stmt_554/forx_xbodyx_xi349_forx_xbodyx_xi349_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(347) & convolution3D_CP_1767_elements(350);
      gj_convolution3D_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  merge  fork  transition  place  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	344 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352: 	354 
    -- CP-element group 352:  members (2) 
      -- CP-element group 352: 	 branch_block_stmt_554/merge_stmt_1563_PhiReqMerge
      -- CP-element group 352: 	 branch_block_stmt_554/merge_stmt_1563_PhiAck/$entry
      -- 
    convolution3D_CP_1767_elements(352) <= OrReduce(convolution3D_CP_1767_elements(344) & convolution3D_CP_1767_elements(351));
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	355 
    -- CP-element group 353:  members (1) 
      -- CP-element group 353: 	 branch_block_stmt_554/merge_stmt_1563_PhiAck/phi_stmt_1564_ack
      -- 
    phi_stmt_1564_ack_4533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1564_ack_0, ack => convolution3D_CP_1767_elements(353)); -- 
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	352 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	355 
    -- CP-element group 354:  members (1) 
      -- CP-element group 354: 	 branch_block_stmt_554/merge_stmt_1563_PhiAck/phi_stmt_1571_ack
      -- 
    phi_stmt_1571_ack_4534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1571_ack_0, ack => convolution3D_CP_1767_elements(354)); -- 
    -- CP-element group 355:  join  fork  transition  place  output  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	353 
    -- CP-element group 355: 	354 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	217 
    -- CP-element group 355: 	218 
    -- CP-element group 355: 	216 
    -- CP-element group 355: 	213 
    -- CP-element group 355:  members (16) 
      -- CP-element group 355: 	 branch_block_stmt_554/merge_stmt_1563__exit__
      -- CP-element group 355: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617__entry__
      -- CP-element group 355: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1596_update_start_
      -- CP-element group 355: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/RPIPE_maxpool_input_pipe_1592_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/RPIPE_maxpool_input_pipe_1592_Sample/rr
      -- CP-element group 355: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/RPIPE_maxpool_input_pipe_1592_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/$entry
      -- CP-element group 355: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1611_Update/cr
      -- CP-element group 355: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1611_Update/$entry
      -- CP-element group 355: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1611_Sample/rr
      -- CP-element group 355: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1611_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1611_update_start_
      -- CP-element group 355: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1611_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1596_Update/cr
      -- CP-element group 355: 	 branch_block_stmt_554/assign_stmt_1584_to_assign_stmt_1617/type_cast_1596_Update/$entry
      -- CP-element group 355: 	 branch_block_stmt_554/merge_stmt_1563_PhiAck/$exit
      -- 
    rr_3508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(355), ack => RPIPE_maxpool_input_pipe_1592_inst_req_0); -- 
    cr_3541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(355), ack => type_cast_1611_inst_req_1); -- 
    rr_3536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(355), ack => type_cast_1611_inst_req_0); -- 
    cr_3527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(355), ack => type_cast_1596_inst_req_1); -- 
    convolution3D_cp_element_group_355: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_355"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(353) & convolution3D_CP_1767_elements(354);
      gj_convolution3D_cp_element_group_355 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(355), clk => clk, reset => reset); --
    end block;
    -- CP-element group 356:  transition  input  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	221 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	358 
    -- CP-element group 356:  members (2) 
      -- CP-element group 356: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1628/SplitProtocol/Sample/$exit
      -- CP-element group 356: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1628/SplitProtocol/Sample/ra
      -- 
    ra_4558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1628_inst_ack_0, ack => convolution3D_CP_1767_elements(356)); -- 
    -- CP-element group 357:  transition  input  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	221 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (2) 
      -- CP-element group 357: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1628/SplitProtocol/Update/ca
      -- CP-element group 357: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1628/SplitProtocol/Update/$exit
      -- 
    ca_4563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1628_inst_ack_1, ack => convolution3D_CP_1767_elements(357)); -- 
    -- CP-element group 358:  join  transition  place  output  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	356 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (8) 
      -- CP-element group 358: 	 branch_block_stmt_554/merge_stmt_1624_PhiReqMerge
      -- CP-element group 358: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1628/$exit
      -- CP-element group 358: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/type_cast_1628/SplitProtocol/$exit
      -- CP-element group 358: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/phi_stmt_1625/phi_stmt_1625_sources/$exit
      -- CP-element group 358: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/phi_stmt_1625/$exit
      -- CP-element group 358: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/$exit
      -- CP-element group 358: 	 branch_block_stmt_554/merge_stmt_1624_PhiAck/$entry
      -- CP-element group 358: 	 branch_block_stmt_554/forx_xbodyx_xi349_getRemainingElementsx_xexit357_PhiReq/phi_stmt_1625/phi_stmt_1625_req
      -- 
    phi_stmt_1625_req_4564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1625_req_4564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(358), ack => phi_stmt_1625_req_0); -- 
    convolution3D_cp_element_group_358: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_358"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(356) & convolution3D_CP_1767_elements(357);
      gj_convolution3D_cp_element_group_358 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(358), clk => clk, reset => reset); --
    end block;
    -- CP-element group 359:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	222 
    -- CP-element group 359: 	223 
    -- CP-element group 359: 	225 
    -- CP-element group 359: 	227 
    -- CP-element group 359:  members (29) 
      -- CP-element group 359: 	 branch_block_stmt_554/merge_stmt_1624__exit__
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663__entry__
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_index_scale_1/scale_rename_ack
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_final_index_sum_regn_update_start
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_final_index_sum_regn_Sample/$entry
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_final_index_sum_regn_Sample/req
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_index_scale_1/scale_rename_req
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_index_scale_1/$exit
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Update/word_access_complete/word_0/cr
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_index_scale_1/$entry
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_index_resize_1/index_resize_ack
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Update/word_access_complete/word_0/$entry
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_index_resize_1/index_resize_req
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_index_resize_1/$exit
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_index_resize_1/$entry
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_index_computed_1
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Update/word_access_complete/$entry
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_index_scaled_1
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_index_resized_1
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_final_index_sum_regn_Update/req
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/addr_of_1658_update_start_
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/array_obj_ref_1657_final_index_sum_regn_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/$entry
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/ptr_deref_1661_update_start_
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/addr_of_1658_complete/req
      -- CP-element group 359: 	 branch_block_stmt_554/assign_stmt_1635_to_assign_stmt_1663/addr_of_1658_complete/$entry
      -- CP-element group 359: 	 branch_block_stmt_554/merge_stmt_1624_PhiAck/phi_stmt_1625_ack
      -- CP-element group 359: 	 branch_block_stmt_554/merge_stmt_1624_PhiAck/$exit
      -- 
    phi_stmt_1625_ack_4569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1625_ack_0, ack => convolution3D_CP_1767_elements(359)); -- 
    req_3589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(359), ack => array_obj_ref_1657_index_offset_req_0); -- 
    cr_3659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(359), ack => ptr_deref_1661_store_0_req_1); -- 
    req_3594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(359), ack => array_obj_ref_1657_index_offset_req_1); -- 
    req_3609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(359), ack => addr_of_1658_final_reg_req_1); -- 
    -- CP-element group 360:  merge  fork  transition  place  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	209 
    -- CP-element group 360: 	228 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	229 
    -- CP-element group 360: 	230 
    -- CP-element group 360:  members (13) 
      -- CP-element group 360: 	 branch_block_stmt_554/merge_stmt_1665__exit__
      -- CP-element group 360: 	 branch_block_stmt_554/call_stmt_1668__entry__
      -- CP-element group 360: 	 branch_block_stmt_554/call_stmt_1668/call_stmt_1668_Sample/$entry
      -- CP-element group 360: 	 branch_block_stmt_554/call_stmt_1668/call_stmt_1668_Sample/crr
      -- CP-element group 360: 	 branch_block_stmt_554/merge_stmt_1665_PhiReqMerge
      -- CP-element group 360: 	 branch_block_stmt_554/call_stmt_1668/call_stmt_1668_Update/$entry
      -- CP-element group 360: 	 branch_block_stmt_554/call_stmt_1668/call_stmt_1668_update_start_
      -- CP-element group 360: 	 branch_block_stmt_554/call_stmt_1668/call_stmt_1668_sample_start_
      -- CP-element group 360: 	 branch_block_stmt_554/call_stmt_1668/$entry
      -- CP-element group 360: 	 branch_block_stmt_554/call_stmt_1668/call_stmt_1668_Update/ccr
      -- CP-element group 360: 	 branch_block_stmt_554/merge_stmt_1665_PhiAck/dummy
      -- CP-element group 360: 	 branch_block_stmt_554/merge_stmt_1665_PhiAck/$exit
      -- CP-element group 360: 	 branch_block_stmt_554/merge_stmt_1665_PhiAck/$entry
      -- 
    crr_3671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(360), ack => call_stmt_1668_call_req_0); -- 
    ccr_3676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(360), ack => call_stmt_1668_call_req_1); -- 
    convolution3D_CP_1767_elements(360) <= OrReduce(convolution3D_CP_1767_elements(209) & convolution3D_CP_1767_elements(228));
    -- CP-element group 361:  transition  output  delay-element  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	239 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	365 
    -- CP-element group 361:  members (5) 
      -- CP-element group 361: 	 branch_block_stmt_554/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_req
      -- CP-element group 361: 	 branch_block_stmt_554/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_sources/type_cast_1716_konst_delay_trans
      -- CP-element group 361: 	 branch_block_stmt_554/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_sources/$exit
      -- CP-element group 361: 	 branch_block_stmt_554/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1710/$exit
      -- CP-element group 361: 	 branch_block_stmt_554/ifx_xend227_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_1710_req_4591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1710_req_4591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(361), ack => phi_stmt_1710_req_1); -- 
    -- Element group convolution3D_CP_1767_elements(361) is a control-delay.
    cp_element_361_delay: control_delay_element  generic map(name => " 361_delay", delay_value => 1)  port map(req => convolution3D_CP_1767_elements(239), ack => convolution3D_CP_1767_elements(361), clk => clk, reset =>reset);
    -- CP-element group 362:  transition  input  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	250 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	364 
    -- CP-element group 362:  members (2) 
      -- CP-element group 362: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_sources/type_cast_1713/SplitProtocol/Sample/ra
      -- CP-element group 362: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_sources/type_cast_1713/SplitProtocol/Sample/$exit
      -- 
    ra_4611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1713_inst_ack_0, ack => convolution3D_CP_1767_elements(362)); -- 
    -- CP-element group 363:  transition  input  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	250 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (2) 
      -- CP-element group 363: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_sources/type_cast_1713/SplitProtocol/Update/ca
      -- CP-element group 363: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_sources/type_cast_1713/SplitProtocol/Update/$exit
      -- 
    ca_4616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1713_inst_ack_1, ack => convolution3D_CP_1767_elements(363)); -- 
    -- CP-element group 364:  join  transition  output  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	362 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (6) 
      -- CP-element group 364: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_req
      -- CP-element group 364: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_sources/type_cast_1713/SplitProtocol/$exit
      -- CP-element group 364: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_sources/type_cast_1713/$exit
      -- CP-element group 364: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1710/phi_stmt_1710_sources/$exit
      -- CP-element group 364: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1710/$exit
      -- CP-element group 364: 	 branch_block_stmt_554/whilex_xbody_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_1710_req_4617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1710_req_4617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(364), ack => phi_stmt_1710_req_0); -- 
    convolution3D_cp_element_group_364: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_364"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1767_elements(362) & convolution3D_CP_1767_elements(363);
      gj_convolution3D_cp_element_group_364 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1767_elements(364), clk => clk, reset => reset); --
    end block;
    -- CP-element group 365:  merge  transition  place  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	361 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (2) 
      -- CP-element group 365: 	 branch_block_stmt_554/merge_stmt_1709_PhiReqMerge
      -- CP-element group 365: 	 branch_block_stmt_554/merge_stmt_1709_PhiAck/$entry
      -- 
    convolution3D_CP_1767_elements(365) <= OrReduce(convolution3D_CP_1767_elements(361) & convolution3D_CP_1767_elements(364));
    -- CP-element group 366:  fork  transition  place  input  output  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	244 
    -- CP-element group 366: 	245 
    -- CP-element group 366: 	246 
    -- CP-element group 366: 	240 
    -- CP-element group 366: 	247 
    -- CP-element group 366:  members (20) 
      -- CP-element group 366: 	 branch_block_stmt_554/merge_stmt_1709__exit__
      -- CP-element group 366: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752__entry__
      -- CP-element group 366: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1723_Sample/req
      -- CP-element group 366: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1741_Update/ccr
      -- CP-element group 366: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1723_Sample/$entry
      -- CP-element group 366: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1741_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1741_Sample/crr
      -- CP-element group 366: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1741_Sample/$entry
      -- CP-element group 366: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1741_update_start_
      -- CP-element group 366: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1741_sample_start_
      -- CP-element group 366: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1737_Update/ccr
      -- CP-element group 366: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1737_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1737_Sample/crr
      -- CP-element group 366: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1737_Sample/$entry
      -- CP-element group 366: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/WPIPE_num_out_pipe_1723_sample_start_
      -- CP-element group 366: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/$entry
      -- CP-element group 366: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1737_update_start_
      -- CP-element group 366: 	 branch_block_stmt_554/assign_stmt_1722_to_assign_stmt_1752/call_stmt_1737_sample_start_
      -- CP-element group 366: 	 branch_block_stmt_554/merge_stmt_1709_PhiAck/phi_stmt_1710_ack
      -- CP-element group 366: 	 branch_block_stmt_554/merge_stmt_1709_PhiAck/$exit
      -- 
    phi_stmt_1710_ack_4622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1710_ack_0, ack => convolution3D_CP_1767_elements(366)); -- 
    req_3747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(366), ack => WPIPE_num_out_pipe_1723_inst_req_0); -- 
    ccr_3794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(366), ack => call_stmt_1741_call_req_1); -- 
    crr_3789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(366), ack => call_stmt_1741_call_req_0); -- 
    ccr_3780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(366), ack => call_stmt_1737_call_req_1); -- 
    crr_3775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1767_elements(366), ack => call_stmt_1737_call_req_0); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i64_i64_1053_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_1240_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_1514_wire : std_logic_vector(63 downto 0);
    signal Bx_xnot_1170 : std_logic_vector(63 downto 0);
    signal R_indvar395_1336_resized : std_logic_vector(13 downto 0);
    signal R_indvar395_1336_scaled : std_logic_vector(13 downto 0);
    signal R_indvar409_875_resized : std_logic_vector(13 downto 0);
    signal R_indvar409_875_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1191_resized : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1191_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1656_resized : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1656_scaled : std_logic_vector(13 downto 0);
    signal add102_921 : std_logic_vector(63 downto 0);
    signal add108_939 : std_logic_vector(63 downto 0);
    signal add114_957 : std_logic_vector(63 downto 0);
    signal add120_975 : std_logic_vector(63 downto 0);
    signal add1216x_xi354_1641 : std_logic_vector(63 downto 0);
    signal add1216x_xi_1176 : std_logic_vector(63 downto 0);
    signal add126_993 : std_logic_vector(63 downto 0);
    signal add132_1011 : std_logic_vector(63 downto 0);
    signal add13_605 : std_logic_vector(15 downto 0);
    signal add171_1364 : std_logic_vector(63 downto 0);
    signal add177_1382 : std_logic_vector(63 downto 0);
    signal add183_1400 : std_logic_vector(63 downto 0);
    signal add189_1418 : std_logic_vector(63 downto 0);
    signal add195_1436 : std_logic_vector(63 downto 0);
    signal add201_1454 : std_logic_vector(63 downto 0);
    signal add207_1472 : std_logic_vector(63 downto 0);
    signal add23_630 : std_logic_vector(15 downto 0);
    signal add33_655 : std_logic_vector(15 downto 0);
    signal add43_680 : std_logic_vector(15 downto 0);
    signal add53_705 : std_logic_vector(15 downto 0);
    signal add63_730 : std_logic_vector(63 downto 0);
    signal add73_755 : std_logic_vector(15 downto 0);
    signal add96_903 : std_logic_vector(63 downto 0);
    signal add_580 : std_logic_vector(31 downto 0);
    signal addx_xi345_1602 : std_logic_vector(63 downto 0);
    signal addx_xi_1137 : std_logic_vector(63 downto 0);
    signal and217_1532 : std_logic_vector(63 downto 0);
    signal and_1071 : std_logic_vector(63 downto 0);
    signal array_obj_ref_1192_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1192_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1192_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1192_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1192_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1192_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1337_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1337_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1337_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1337_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1337_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1337_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1657_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1657_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1657_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1657_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1657_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1657_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_876_root_address : std_logic_vector(13 downto 0);
    signal arrayidx143_1194 : std_logic_vector(31 downto 0);
    signal arrayidx211_1339 : std_logic_vector(31 downto 0);
    signal arrayidx226_1659 : std_logic_vector(31 downto 0);
    signal arrayidx_878 : std_logic_vector(31 downto 0);
    signal call105_930 : std_logic_vector(7 downto 0);
    signal call111_948 : std_logic_vector(7 downto 0);
    signal call117_966 : std_logic_vector(7 downto 0);
    signal call11_596 : std_logic_vector(7 downto 0);
    signal call123_984 : std_logic_vector(7 downto 0);
    signal call129_1002 : std_logic_vector(7 downto 0);
    signal call164_1342 : std_logic_vector(7 downto 0);
    signal call168_1355 : std_logic_vector(7 downto 0);
    signal call16_608 : std_logic_vector(7 downto 0);
    signal call174_1373 : std_logic_vector(7 downto 0);
    signal call180_1391 : std_logic_vector(7 downto 0);
    signal call186_1409 : std_logic_vector(7 downto 0);
    signal call192_1427 : std_logic_vector(7 downto 0);
    signal call198_1445 : std_logic_vector(7 downto 0);
    signal call204_1463 : std_logic_vector(7 downto 0);
    signal call21_621 : std_logic_vector(7 downto 0);
    signal call229_1668 : std_logic_vector(63 downto 0);
    signal call267_1767 : std_logic_vector(7 downto 0);
    signal call269_1770 : std_logic_vector(63 downto 0);
    signal call26_633 : std_logic_vector(7 downto 0);
    signal call2_571 : std_logic_vector(7 downto 0);
    signal call31_646 : std_logic_vector(7 downto 0);
    signal call36_658 : std_logic_vector(7 downto 0);
    signal call41_671 : std_logic_vector(7 downto 0);
    signal call46_683 : std_logic_vector(7 downto 0);
    signal call51_696 : std_logic_vector(7 downto 0);
    signal call56_708 : std_logic_vector(7 downto 0);
    signal call61_721 : std_logic_vector(7 downto 0);
    signal call66_733 : std_logic_vector(7 downto 0);
    signal call6_583 : std_logic_vector(7 downto 0);
    signal call71_746 : std_logic_vector(7 downto 0);
    signal call89_881 : std_logic_vector(7 downto 0);
    signal call93_894 : std_logic_vector(7 downto 0);
    signal call99_912 : std_logic_vector(7 downto 0);
    signal call_558 : std_logic_vector(7 downto 0);
    signal callx_xi343_1593 : std_logic_vector(7 downto 0);
    signal callx_xi_1128 : std_logic_vector(7 downto 0);
    signal cmp161363_1248 : std_logic_vector(0 downto 0);
    signal cmp367_785 : std_logic_vector(0 downto 0);
    signal cmpx_xi348_1617 : std_logic_vector(0 downto 0);
    signal cmpx_xi_1152 : std_logic_vector(0 downto 0);
    signal conv101_916 : std_logic_vector(63 downto 0);
    signal conv107_934 : std_logic_vector(63 downto 0);
    signal conv113_952 : std_logic_vector(63 downto 0);
    signal conv119_970 : std_logic_vector(63 downto 0);
    signal conv125_988 : std_logic_vector(63 downto 0);
    signal conv12_600 : std_logic_vector(15 downto 0);
    signal conv131_1006 : std_logic_vector(63 downto 0);
    signal conv145_1204 : std_logic_vector(63 downto 0);
    signal conv147_1208 : std_logic_vector(63 downto 0);
    signal conv153_1212 : std_logic_vector(63 downto 0);
    signal conv155_1242 : std_logic_vector(63 downto 0);
    signal conv165_1346 : std_logic_vector(63 downto 0);
    signal conv170_1359 : std_logic_vector(63 downto 0);
    signal conv176_1377 : std_logic_vector(63 downto 0);
    signal conv182_1395 : std_logic_vector(63 downto 0);
    signal conv188_1413 : std_logic_vector(63 downto 0);
    signal conv194_1431 : std_logic_vector(63 downto 0);
    signal conv19_612 : std_logic_vector(15 downto 0);
    signal conv1_562 : std_logic_vector(31 downto 0);
    signal conv200_1449 : std_logic_vector(63 downto 0);
    signal conv206_1467 : std_logic_vector(63 downto 0);
    signal conv22_625 : std_logic_vector(15 downto 0);
    signal conv230_1764 : std_logic_vector(63 downto 0);
    signal conv251_1734 : std_logic_vector(63 downto 0);
    signal conv270_1775 : std_logic_vector(63 downto 0);
    signal conv277_1784 : std_logic_vector(7 downto 0);
    signal conv283_1794 : std_logic_vector(7 downto 0);
    signal conv289_1804 : std_logic_vector(7 downto 0);
    signal conv295_1814 : std_logic_vector(7 downto 0);
    signal conv29_637 : std_logic_vector(15 downto 0);
    signal conv2x_xi338_1555 : std_logic_vector(31 downto 0);
    signal conv2x_xi_1090 : std_logic_vector(31 downto 0);
    signal conv301_1824 : std_logic_vector(7 downto 0);
    signal conv307_1834 : std_logic_vector(7 downto 0);
    signal conv313_1844 : std_logic_vector(7 downto 0);
    signal conv319_1854 : std_logic_vector(7 downto 0);
    signal conv32_650 : std_logic_vector(15 downto 0);
    signal conv39_662 : std_logic_vector(15 downto 0);
    signal conv3_575 : std_logic_vector(31 downto 0);
    signal conv42_675 : std_logic_vector(15 downto 0);
    signal conv49_687 : std_logic_vector(15 downto 0);
    signal conv52_700 : std_logic_vector(15 downto 0);
    signal conv59_712 : std_logic_vector(63 downto 0);
    signal conv5x_xi344_1597 : std_logic_vector(63 downto 0);
    signal conv5x_xi_1132 : std_logic_vector(63 downto 0);
    signal conv62_725 : std_logic_vector(63 downto 0);
    signal conv69_737 : std_logic_vector(15 downto 0);
    signal conv72_750 : std_logic_vector(15 downto 0);
    signal conv79_759 : std_logic_vector(31 downto 0);
    signal conv81_763 : std_logic_vector(31 downto 0);
    signal conv83_779 : std_logic_vector(63 downto 0);
    signal conv90_885 : std_logic_vector(63 downto 0);
    signal conv95_898 : std_logic_vector(63 downto 0);
    signal conv9_587 : std_logic_vector(15 downto 0);
    signal convx_xi347_1612 : std_logic_vector(31 downto 0);
    signal convx_xi_1147 : std_logic_vector(31 downto 0);
    signal elementx_x021x_xi342_1571 : std_logic_vector(63 downto 0);
    signal elementx_x021x_xi_1106 : std_logic_vector(63 downto 0);
    signal exitcond28_1026 : std_logic_vector(0 downto 0);
    signal exitcond5_1752 : std_logic_vector(0 downto 0);
    signal exitcond_1487 : std_logic_vector(0 downto 0);
    signal iNsTr_35_1125 : std_logic_vector(15 downto 0);
    signal iNsTr_55_1551 : std_logic_vector(63 downto 0);
    signal iNsTr_67_1590 : std_logic_vector(15 downto 0);
    signal iNsTr_90_1635 : std_logic_vector(63 downto 0);
    signal indvar395_1325 : std_logic_vector(63 downto 0);
    signal indvar409_864 : std_logic_vector(63 downto 0);
    signal indvar_1710 : std_logic_vector(63 downto 0);
    signal indvarx_xnext396_1482 : std_logic_vector(63 downto 0);
    signal indvarx_xnext410_1021 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1747 : std_logic_vector(63 downto 0);
    signal ix_x0x_xlcssa_1058 : std_logic_vector(63 downto 0);
    signal ix_x1x_xlcssa_1519 : std_logic_vector(63 downto 0);
    signal mul148_1217 : std_logic_vector(63 downto 0);
    signal mul151_1222 : std_logic_vector(63 downto 0);
    signal mul154_1227 : std_logic_vector(63 downto 0);
    signal mul250_1722 : std_logic_vector(63 downto 0);
    signal mul82_773 : std_logic_vector(31 downto 0);
    signal mul_768 : std_logic_vector(31 downto 0);
    signal nx_x022x_xi341_1564 : std_logic_vector(15 downto 0);
    signal nx_x022x_xi_1099 : std_logic_vector(15 downto 0);
    signal phitmp371_1516 : std_logic_vector(63 downto 0);
    signal phitmp_1055 : std_logic_vector(63 downto 0);
    signal ptr_deref_1013_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1013_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1013_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1013_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1013_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1013_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1196_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1196_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1196_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1196_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1196_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1196_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1474_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1474_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1474_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1474_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1474_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1474_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1661_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1661_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1661_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1661_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1661_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1661_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext_1233 : std_logic_vector(63 downto 0);
    signal sh_promx_xi355_1647 : std_logic_vector(63 downto 0);
    signal sh_promx_xi_1182 : std_logic_vector(63 downto 0);
    signal shl104_927 : std_logic_vector(63 downto 0);
    signal shl10_593 : std_logic_vector(15 downto 0);
    signal shl110_945 : std_logic_vector(63 downto 0);
    signal shl116_963 : std_logic_vector(63 downto 0);
    signal shl122_981 : std_logic_vector(63 downto 0);
    signal shl128_999 : std_logic_vector(63 downto 0);
    signal shl14x_xi356_1652 : std_logic_vector(63 downto 0);
    signal shl14x_xi_1187 : std_logic_vector(63 downto 0);
    signal shl167_1352 : std_logic_vector(63 downto 0);
    signal shl173_1370 : std_logic_vector(63 downto 0);
    signal shl179_1388 : std_logic_vector(63 downto 0);
    signal shl185_1406 : std_logic_vector(63 downto 0);
    signal shl191_1424 : std_logic_vector(63 downto 0);
    signal shl197_1442 : std_logic_vector(63 downto 0);
    signal shl203_1460 : std_logic_vector(63 downto 0);
    signal shl20_618 : std_logic_vector(15 downto 0);
    signal shl30_643 : std_logic_vector(15 downto 0);
    signal shl40_668 : std_logic_vector(15 downto 0);
    signal shl50_693 : std_logic_vector(15 downto 0);
    signal shl60_718 : std_logic_vector(63 downto 0);
    signal shl70_743 : std_logic_vector(15 downto 0);
    signal shl8x_xi346_1608 : std_logic_vector(63 downto 0);
    signal shl8x_xi346x_xlcssa_1625 : std_logic_vector(63 downto 0);
    signal shl8x_xi_1143 : std_logic_vector(63 downto 0);
    signal shl8x_xix_xlcssa_1160 : std_logic_vector(63 downto 0);
    signal shl92_891 : std_logic_vector(63 downto 0);
    signal shl98_909 : std_logic_vector(63 downto 0);
    signal shl_568 : std_logic_vector(31 downto 0);
    signal shlx_xi339_1561 : std_logic_vector(31 downto 0);
    signal shlx_xi_1096 : std_logic_vector(31 downto 0);
    signal shr280_1790 : std_logic_vector(63 downto 0);
    signal shr286_1800 : std_logic_vector(63 downto 0);
    signal shr292_1810 : std_logic_vector(63 downto 0);
    signal shr298_1820 : std_logic_vector(63 downto 0);
    signal shr304_1830 : std_logic_vector(63 downto 0);
    signal shr310_1840 : std_logic_vector(63 downto 0);
    signal shr316_1850 : std_logic_vector(63 downto 0);
    signal sub_1780 : std_logic_vector(63 downto 0);
    signal tmp10_1276 : std_logic_vector(63 downto 0);
    signal tmp11_1280 : std_logic_vector(63 downto 0);
    signal tmp12_1285 : std_logic_vector(63 downto 0);
    signal tmp13_1289 : std_logic_vector(63 downto 0);
    signal tmp14_1294 : std_logic_vector(63 downto 0);
    signal tmp15_1298 : std_logic_vector(31 downto 0);
    signal tmp16_1303 : std_logic_vector(63 downto 0);
    signal tmp17_1309 : std_logic_vector(63 downto 0);
    signal tmp18_1315 : std_logic_vector(0 downto 0);
    signal tmp20_823 : std_logic_vector(31 downto 0);
    signal tmp21_828 : std_logic_vector(31 downto 0);
    signal tmp22_832 : std_logic_vector(31 downto 0);
    signal tmp23_837 : std_logic_vector(31 downto 0);
    signal tmp24_842 : std_logic_vector(63 downto 0);
    signal tmp25_848 : std_logic_vector(63 downto 0);
    signal tmp26_854 : std_logic_vector(0 downto 0);
    signal tmp372_1584 : std_logic_vector(15 downto 0);
    signal tmp373_1683 : std_logic_vector(15 downto 0);
    signal tmp377_1688 : std_logic_vector(15 downto 0);
    signal tmp390_1261 : std_logic_vector(63 downto 0);
    signal tmp391_1267 : std_logic_vector(0 downto 0);
    signal tmp392_1507 : std_logic_vector(63 downto 0);
    signal tmp399_797 : std_logic_vector(31 downto 0);
    signal tmp3_1692 : std_logic_vector(63 downto 0);
    signal tmp401_802 : std_logic_vector(31 downto 0);
    signal tmp402_807 : std_logic_vector(63 downto 0);
    signal tmp403_813 : std_logic_vector(63 downto 0);
    signal tmp404_819 : std_logic_vector(0 downto 0);
    signal tmp406_1046 : std_logic_vector(63 downto 0);
    signal tmp4_1698 : std_logic_vector(63 downto 0);
    signal tmp6_1702 : std_logic_vector(63 downto 0);
    signal tmp7_1707 : std_logic_vector(63 downto 0);
    signal tmp9_1271 : std_logic_vector(63 downto 0);
    signal tmp_1119 : std_logic_vector(15 downto 0);
    signal tobool218_1538 : std_logic_vector(0 downto 0);
    signal tobool_1077 : std_logic_vector(0 downto 0);
    signal type_cast_1019_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1038_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1044_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1049_wire : std_logic_vector(63 downto 0);
    signal type_cast_1052_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1061_wire : std_logic_vector(63 downto 0);
    signal type_cast_1064_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1069_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1075_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1088_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1094_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1103_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1105_wire : std_logic_vector(15 downto 0);
    signal type_cast_1110_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1112_wire : std_logic_vector(63 downto 0);
    signal type_cast_1117_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1123_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1141_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1163_wire : std_logic_vector(63 downto 0);
    signal type_cast_1168_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1174_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1180_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1231_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1236_wire : std_logic_vector(63 downto 0);
    signal type_cast_1239_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1246_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1259_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1265_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1301_wire : std_logic_vector(63 downto 0);
    signal type_cast_1307_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1313_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1320_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1329_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1331_wire : std_logic_vector(63 downto 0);
    signal type_cast_1350_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1368_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1386_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1404_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1422_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1440_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1458_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1480_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1499_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1505_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1510_wire : std_logic_vector(63 downto 0);
    signal type_cast_1513_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1522_wire : std_logic_vector(63 downto 0);
    signal type_cast_1525_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1530_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1536_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1549_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1559_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1568_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1570_wire : std_logic_vector(15 downto 0);
    signal type_cast_1575_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1577_wire : std_logic_vector(63 downto 0);
    signal type_cast_1582_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1588_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1606_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1628_wire : std_logic_vector(63 downto 0);
    signal type_cast_1633_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1639_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1645_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1672_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1676_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1681_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1696_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1713_wire : std_logic_vector(63 downto 0);
    signal type_cast_1716_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1732_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1745_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1762_wire : std_logic_vector(63 downto 0);
    signal type_cast_1773_wire : std_logic_vector(63 downto 0);
    signal type_cast_1788_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1798_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1808_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1818_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1828_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1838_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1848_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_566_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_591_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_616_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_641_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_666_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_691_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_716_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_741_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_777_wire : std_logic_vector(63 downto 0);
    signal type_cast_783_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_805_wire : std_logic_vector(63 downto 0);
    signal type_cast_811_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_817_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_840_wire : std_logic_vector(63 downto 0);
    signal type_cast_846_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_852_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_859_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_868_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_870_wire : std_logic_vector(63 downto 0);
    signal type_cast_889_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_907_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_925_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_943_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_961_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_979_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_997_wire_constant : std_logic_vector(63 downto 0);
    signal umax19_1322 : std_logic_vector(63 downto 0);
    signal umax27_861 : std_logic_vector(63 downto 0);
    signal umax405_1040 : std_logic_vector(63 downto 0);
    signal umax_1501 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1192_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1192_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1192_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1192_resized_base_address <= "00000000000000";
    array_obj_ref_1337_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1337_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1337_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1337_resized_base_address <= "00000000000000";
    array_obj_ref_1657_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1657_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1657_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1657_resized_base_address <= "00000000000000";
    array_obj_ref_876_constant_part_of_offset <= "00000000000000";
    array_obj_ref_876_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_876_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_876_resized_base_address <= "00000000000000";
    ptr_deref_1013_word_offset_0 <= "00000000000000";
    ptr_deref_1196_word_offset_0 <= "00000000000000";
    ptr_deref_1474_word_offset_0 <= "00000000000000";
    ptr_deref_1661_word_offset_0 <= "00000000000000";
    type_cast_1019_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1038_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1044_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1052_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1064_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1069_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1075_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1088_wire_constant <= "00000000000000000000000000000001";
    type_cast_1094_wire_constant <= "00000000000000000000000000000110";
    type_cast_1103_wire_constant <= "0000000000000000";
    type_cast_1110_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1117_wire_constant <= "0000000000000001";
    type_cast_1123_wire_constant <= "0000000000000001";
    type_cast_1141_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1168_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1174_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1180_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1231_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1239_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1246_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1259_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1265_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1307_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1313_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1320_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1329_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1350_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1368_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1386_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1404_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1422_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1440_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1458_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1480_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1499_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1505_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1513_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1525_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1530_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1536_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1549_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1559_wire_constant <= "00000000000000000000000000000110";
    type_cast_1568_wire_constant <= "0000000000000000";
    type_cast_1575_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1582_wire_constant <= "0000000000000001";
    type_cast_1588_wire_constant <= "0000000000000001";
    type_cast_1606_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1633_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1639_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1645_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1672_wire_constant <= "11001000";
    type_cast_1676_wire_constant <= "11001000";
    type_cast_1681_wire_constant <= "1111111111111111";
    type_cast_1696_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1716_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1732_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111111";
    type_cast_1745_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1788_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1798_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1808_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1818_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1828_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1838_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1848_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_566_wire_constant <= "00000000000000000000000000001000";
    type_cast_591_wire_constant <= "0000000000001000";
    type_cast_616_wire_constant <= "0000000000001000";
    type_cast_641_wire_constant <= "0000000000001000";
    type_cast_666_wire_constant <= "0000000000001000";
    type_cast_691_wire_constant <= "0000000000001000";
    type_cast_716_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_741_wire_constant <= "0000000000001000";
    type_cast_783_wire_constant <= "00000000000000000000000000000011";
    type_cast_811_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_817_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_846_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_852_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_859_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_868_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_889_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_907_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_925_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_943_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_961_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_979_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_997_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    phi_stmt_1058: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1061_wire & type_cast_1064_wire_constant;
      req <= phi_stmt_1058_req_0 & phi_stmt_1058_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1058",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1058_ack_0,
          idata => idata,
          odata => ix_x0x_xlcssa_1058,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1058
    phi_stmt_1099: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1103_wire_constant & type_cast_1105_wire;
      req <= phi_stmt_1099_req_0 & phi_stmt_1099_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1099",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1099_ack_0,
          idata => idata,
          odata => nx_x022x_xi_1099,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1099
    phi_stmt_1106: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1110_wire_constant & type_cast_1112_wire;
      req <= phi_stmt_1106_req_0 & phi_stmt_1106_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1106",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1106_ack_0,
          idata => idata,
          odata => elementx_x021x_xi_1106,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1106
    phi_stmt_1160: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1163_wire;
      req(0) <= phi_stmt_1160_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1160",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1160_ack_0,
          idata => idata,
          odata => shl8x_xix_xlcssa_1160,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1160
    phi_stmt_1325: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1329_wire_constant & type_cast_1331_wire;
      req <= phi_stmt_1325_req_0 & phi_stmt_1325_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1325",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1325_ack_0,
          idata => idata,
          odata => indvar395_1325,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1325
    phi_stmt_1519: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1522_wire & type_cast_1525_wire_constant;
      req <= phi_stmt_1519_req_0 & phi_stmt_1519_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1519",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1519_ack_0,
          idata => idata,
          odata => ix_x1x_xlcssa_1519,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1519
    phi_stmt_1564: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1568_wire_constant & type_cast_1570_wire;
      req <= phi_stmt_1564_req_0 & phi_stmt_1564_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1564",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1564_ack_0,
          idata => idata,
          odata => nx_x022x_xi341_1564,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1564
    phi_stmt_1571: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1575_wire_constant & type_cast_1577_wire;
      req <= phi_stmt_1571_req_0 & phi_stmt_1571_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1571",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1571_ack_0,
          idata => idata,
          odata => elementx_x021x_xi342_1571,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1571
    phi_stmt_1625: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1628_wire;
      req(0) <= phi_stmt_1625_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1625",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1625_ack_0,
          idata => idata,
          odata => shl8x_xi346x_xlcssa_1625,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1625
    phi_stmt_1710: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1713_wire & type_cast_1716_wire_constant;
      req <= phi_stmt_1710_req_0 & phi_stmt_1710_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1710",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1710_ack_0,
          idata => idata,
          odata => indvar_1710,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1710
    phi_stmt_864: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_868_wire_constant & type_cast_870_wire;
      req <= phi_stmt_864_req_0 & phi_stmt_864_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_864",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_864_ack_0,
          idata => idata,
          odata => indvar409_864,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_864
    -- flow-through select operator MUX_1039_inst
    umax405_1040 <= tmp403_813 when (tmp404_819(0) /=  '0') else type_cast_1038_wire_constant;
    -- flow-through select operator MUX_1321_inst
    umax19_1322 <= tmp17_1309 when (tmp18_1315(0) /=  '0') else type_cast_1320_wire_constant;
    -- flow-through select operator MUX_1500_inst
    umax_1501 <= tmp390_1261 when (tmp391_1267(0) /=  '0') else type_cast_1499_wire_constant;
    -- flow-through select operator MUX_860_inst
    umax27_861 <= tmp25_848 when (tmp26_854(0) /=  '0') else type_cast_859_wire_constant;
    addr_of_1193_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1193_final_reg_req_0;
      addr_of_1193_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1193_final_reg_req_1;
      addr_of_1193_final_reg_ack_1<= rack(0);
      addr_of_1193_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1193_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1192_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx143_1194,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1338_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1338_final_reg_req_0;
      addr_of_1338_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1338_final_reg_req_1;
      addr_of_1338_final_reg_ack_1<= rack(0);
      addr_of_1338_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1338_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1337_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx211_1339,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1658_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1658_final_reg_req_0;
      addr_of_1658_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1658_final_reg_req_1;
      addr_of_1658_final_reg_ack_1<= rack(0);
      addr_of_1658_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1658_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1657_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx226_1659,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_877_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_877_final_reg_req_0;
      addr_of_877_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_877_final_reg_req_1;
      addr_of_877_final_reg_ack_1<= rack(0);
      addr_of_877_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_877_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_876_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_878,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1005_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1005_inst_req_0;
      type_cast_1005_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1005_inst_req_1;
      type_cast_1005_inst_ack_1<= rack(0);
      type_cast_1005_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1005_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call129_1002,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_1006,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1049_inst
    process(tmp406_1046) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp406_1046(63 downto 0);
      type_cast_1049_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1054_inst
    process(ASHR_i64_i64_1053_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1053_wire(63 downto 0);
      phitmp_1055 <= tmp_var; -- 
    end process;
    type_cast_1061_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1061_inst_req_0;
      type_cast_1061_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1061_inst_req_1;
      type_cast_1061_inst_ack_1<= rack(0);
      type_cast_1061_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1061_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp_1055,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1061_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1105_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1105_inst_req_0;
      type_cast_1105_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1105_inst_req_1;
      type_cast_1105_inst_ack_1<= rack(0);
      type_cast_1105_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1105_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_35_1125,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1105_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1112_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1112_inst_req_0;
      type_cast_1112_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1112_inst_req_1;
      type_cast_1112_inst_ack_1<= rack(0);
      type_cast_1112_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1112_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi_1143,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1112_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1131_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1131_inst_req_0;
      type_cast_1131_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1131_inst_req_1;
      type_cast_1131_inst_ack_1<= rack(0);
      type_cast_1131_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1131_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi_1128,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi_1132,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1146_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1146_inst_req_0;
      type_cast_1146_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1146_inst_req_1;
      type_cast_1146_inst_ack_1<= rack(0);
      type_cast_1146_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1146_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_1119,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi_1147,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1163_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1163_inst_req_0;
      type_cast_1163_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1163_inst_req_1;
      type_cast_1163_inst_ack_1<= rack(0);
      type_cast_1163_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1163_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi_1143,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1163_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1203_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1203_inst_req_0;
      type_cast_1203_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1203_inst_req_1;
      type_cast_1203_inst_ack_1<= rack(0);
      type_cast_1203_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1203_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_630,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv145_1204,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1207_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1207_inst_req_0;
      type_cast_1207_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1207_inst_req_1;
      type_cast_1207_inst_ack_1<= rack(0);
      type_cast_1207_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1207_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_755,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_1208,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1211_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1211_inst_req_0;
      type_cast_1211_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1211_inst_req_1;
      type_cast_1211_inst_ack_1<= rack(0);
      type_cast_1211_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1211_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_705,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_1212,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1236_inst
    process(sext_1233) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext_1233(63 downto 0);
      type_cast_1236_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1241_inst
    process(ASHR_i64_i64_1240_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1240_wire(63 downto 0);
      conv155_1242 <= tmp_var; -- 
    end process;
    type_cast_1270_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1270_inst_req_0;
      type_cast_1270_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1270_inst_req_1;
      type_cast_1270_inst_ack_1<= rack(0);
      type_cast_1270_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1270_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_705,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp9_1271,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1279_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1279_inst_req_0;
      type_cast_1279_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1279_inst_req_1;
      type_cast_1279_inst_ack_1<= rack(0);
      type_cast_1279_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1279_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_630,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp11_1280,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1288_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1288_inst_req_0;
      type_cast_1288_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1288_inst_req_1;
      type_cast_1288_inst_ack_1<= rack(0);
      type_cast_1288_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1288_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_755,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp13_1289,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1297_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1297_inst_req_0;
      type_cast_1297_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1297_inst_req_1;
      type_cast_1297_inst_ack_1<= rack(0);
      type_cast_1297_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1297_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp14_1294,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp15_1298,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1302_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1302_inst_req_0;
      type_cast_1302_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1302_inst_req_1;
      type_cast_1302_inst_ack_1<= rack(0);
      type_cast_1302_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1302_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1301_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp16_1303,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1331_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1331_inst_req_0;
      type_cast_1331_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1331_inst_req_1;
      type_cast_1331_inst_ack_1<= rack(0);
      type_cast_1331_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1331_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext396_1482,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1331_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1345_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1345_inst_req_0;
      type_cast_1345_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1345_inst_req_1;
      type_cast_1345_inst_ack_1<= rack(0);
      type_cast_1345_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1345_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call164_1342,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_1346,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1358_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1358_inst_req_0;
      type_cast_1358_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1358_inst_req_1;
      type_cast_1358_inst_ack_1<= rack(0);
      type_cast_1358_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1358_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call168_1355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv170_1359,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1376_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1376_inst_req_0;
      type_cast_1376_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1376_inst_req_1;
      type_cast_1376_inst_ack_1<= rack(0);
      type_cast_1376_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1376_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call174_1373,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv176_1377,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1394_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1394_inst_req_0;
      type_cast_1394_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1394_inst_req_1;
      type_cast_1394_inst_ack_1<= rack(0);
      type_cast_1394_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1394_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call180_1391,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv182_1395,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1412_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1412_inst_req_0;
      type_cast_1412_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1412_inst_req_1;
      type_cast_1412_inst_ack_1<= rack(0);
      type_cast_1412_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1412_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call186_1409,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv188_1413,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1430_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1430_inst_req_0;
      type_cast_1430_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1430_inst_req_1;
      type_cast_1430_inst_ack_1<= rack(0);
      type_cast_1430_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1430_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call192_1427,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv194_1431,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1448_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1448_inst_req_0;
      type_cast_1448_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1448_inst_req_1;
      type_cast_1448_inst_ack_1<= rack(0);
      type_cast_1448_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1448_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call198_1445,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_1449,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1466_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1466_inst_req_0;
      type_cast_1466_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1466_inst_req_1;
      type_cast_1466_inst_ack_1<= rack(0);
      type_cast_1466_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1466_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call204_1463,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv206_1467,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1510_inst
    process(tmp392_1507) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp392_1507(63 downto 0);
      type_cast_1510_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1515_inst
    process(ASHR_i64_i64_1514_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1514_wire(63 downto 0);
      phitmp371_1516 <= tmp_var; -- 
    end process;
    type_cast_1522_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1522_inst_req_0;
      type_cast_1522_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1522_inst_req_1;
      type_cast_1522_inst_ack_1<= rack(0);
      type_cast_1522_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1522_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp371_1516,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1522_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1554_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1554_inst_req_0;
      type_cast_1554_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1554_inst_req_1;
      type_cast_1554_inst_ack_1<= rack(0);
      type_cast_1554_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1554_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_55_1551,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2x_xi338_1555,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1570_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1570_inst_req_0;
      type_cast_1570_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1570_inst_req_1;
      type_cast_1570_inst_ack_1<= rack(0);
      type_cast_1570_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1570_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_67_1590,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1570_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1577_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1577_inst_req_0;
      type_cast_1577_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1577_inst_req_1;
      type_cast_1577_inst_ack_1<= rack(0);
      type_cast_1577_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1577_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi346_1608,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1577_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1596_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1596_inst_req_0;
      type_cast_1596_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1596_inst_req_1;
      type_cast_1596_inst_ack_1<= rack(0);
      type_cast_1596_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1596_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi343_1593,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi344_1597,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1611_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1611_inst_req_0;
      type_cast_1611_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1611_inst_req_1;
      type_cast_1611_inst_ack_1<= rack(0);
      type_cast_1611_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1611_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp372_1584,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi347_1612,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1628_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1628_inst_req_0;
      type_cast_1628_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1628_inst_req_1;
      type_cast_1628_inst_ack_1<= rack(0);
      type_cast_1628_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1628_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi346_1608,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1628_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1691_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1691_inst_req_0;
      type_cast_1691_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1691_inst_req_1;
      type_cast_1691_inst_ack_1<= rack(0);
      type_cast_1691_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1691_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp373_1683,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_1692,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1701_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1701_inst_req_0;
      type_cast_1701_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1701_inst_req_1;
      type_cast_1701_inst_ack_1<= rack(0);
      type_cast_1701_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1701_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp377_1688,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp6_1702,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1713_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1713_inst_req_0;
      type_cast_1713_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1713_inst_req_1;
      type_cast_1713_inst_ack_1<= rack(0);
      type_cast_1713_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1713_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1747,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1713_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1763_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1763_inst_req_0;
      type_cast_1763_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1763_inst_req_1;
      type_cast_1763_inst_ack_1<= rack(0);
      type_cast_1763_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1763_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1762_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv230_1764,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1774_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1774_inst_req_0;
      type_cast_1774_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1774_inst_req_1;
      type_cast_1774_inst_ack_1<= rack(0);
      type_cast_1774_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1774_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1773_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv270_1775,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1783_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1783_inst_req_0;
      type_cast_1783_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1783_inst_req_1;
      type_cast_1783_inst_ack_1<= rack(0);
      type_cast_1783_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1783_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1780,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv277_1784,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1793_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1793_inst_req_0;
      type_cast_1793_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1793_inst_req_1;
      type_cast_1793_inst_ack_1<= rack(0);
      type_cast_1793_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1793_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr280_1790,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv283_1794,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1803_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1803_inst_req_0;
      type_cast_1803_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1803_inst_req_1;
      type_cast_1803_inst_ack_1<= rack(0);
      type_cast_1803_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1803_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr286_1800,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv289_1804,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1813_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1813_inst_req_0;
      type_cast_1813_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1813_inst_req_1;
      type_cast_1813_inst_ack_1<= rack(0);
      type_cast_1813_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1813_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr292_1810,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv295_1814,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1823_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1823_inst_req_0;
      type_cast_1823_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1823_inst_req_1;
      type_cast_1823_inst_ack_1<= rack(0);
      type_cast_1823_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1823_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr298_1820,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv301_1824,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1833_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1833_inst_req_0;
      type_cast_1833_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1833_inst_req_1;
      type_cast_1833_inst_ack_1<= rack(0);
      type_cast_1833_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1833_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr304_1830,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv307_1834,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1843_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1843_inst_req_0;
      type_cast_1843_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1843_inst_req_1;
      type_cast_1843_inst_ack_1<= rack(0);
      type_cast_1843_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1843_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr310_1840,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv313_1844,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1853_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1853_inst_req_0;
      type_cast_1853_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1853_inst_req_1;
      type_cast_1853_inst_ack_1<= rack(0);
      type_cast_1853_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1853_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr316_1850,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv319_1854,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_561_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_561_inst_req_0;
      type_cast_561_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_561_inst_req_1;
      type_cast_561_inst_ack_1<= rack(0);
      type_cast_561_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_561_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_558,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_562,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_574_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_574_inst_req_0;
      type_cast_574_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_574_inst_req_1;
      type_cast_574_inst_ack_1<= rack(0);
      type_cast_574_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_574_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_571,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_575,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_586_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_586_inst_req_0;
      type_cast_586_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_586_inst_req_1;
      type_cast_586_inst_ack_1<= rack(0);
      type_cast_586_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_586_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_583,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_587,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_599_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_599_inst_req_0;
      type_cast_599_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_599_inst_req_1;
      type_cast_599_inst_ack_1<= rack(0);
      type_cast_599_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_599_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_596,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_600,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_611_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_611_inst_req_0;
      type_cast_611_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_611_inst_req_1;
      type_cast_611_inst_ack_1<= rack(0);
      type_cast_611_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_611_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_608,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_612,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_624_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_624_inst_req_0;
      type_cast_624_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_624_inst_req_1;
      type_cast_624_inst_ack_1<= rack(0);
      type_cast_624_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_624_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call21_621,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_625,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_636_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_636_inst_req_0;
      type_cast_636_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_636_inst_req_1;
      type_cast_636_inst_ack_1<= rack(0);
      type_cast_636_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_636_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_633,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_637,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_649_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_649_inst_req_0;
      type_cast_649_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_649_inst_req_1;
      type_cast_649_inst_ack_1<= rack(0);
      type_cast_649_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_649_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_646,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_650,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_661_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_661_inst_req_0;
      type_cast_661_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_661_inst_req_1;
      type_cast_661_inst_ack_1<= rack(0);
      type_cast_661_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_661_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_658,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_662,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_674_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_674_inst_req_0;
      type_cast_674_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_674_inst_req_1;
      type_cast_674_inst_ack_1<= rack(0);
      type_cast_674_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_674_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_671,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_675,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_686_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_686_inst_req_0;
      type_cast_686_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_686_inst_req_1;
      type_cast_686_inst_ack_1<= rack(0);
      type_cast_686_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_686_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_683,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_687,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_699_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_699_inst_req_0;
      type_cast_699_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_699_inst_req_1;
      type_cast_699_inst_ack_1<= rack(0);
      type_cast_699_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_699_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call51_696,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_700,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_711_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_711_inst_req_0;
      type_cast_711_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_711_inst_req_1;
      type_cast_711_inst_ack_1<= rack(0);
      type_cast_711_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_711_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call56_708,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_712,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_724_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_724_inst_req_0;
      type_cast_724_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_724_inst_req_1;
      type_cast_724_inst_ack_1<= rack(0);
      type_cast_724_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_724_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call61_721,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_725,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_736_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_736_inst_req_0;
      type_cast_736_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_736_inst_req_1;
      type_cast_736_inst_ack_1<= rack(0);
      type_cast_736_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_736_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call66_733,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_737,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_749_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_749_inst_req_0;
      type_cast_749_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_749_inst_req_1;
      type_cast_749_inst_ack_1<= rack(0);
      type_cast_749_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_749_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call71_746,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv72_750,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_758_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_758_inst_req_0;
      type_cast_758_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_758_inst_req_1;
      type_cast_758_inst_ack_1<= rack(0);
      type_cast_758_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_758_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_605,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_759,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_762_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_762_inst_req_0;
      type_cast_762_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_762_inst_req_1;
      type_cast_762_inst_ack_1<= rack(0);
      type_cast_762_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_762_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_630,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv81_763,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_778_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_778_inst_req_0;
      type_cast_778_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_778_inst_req_1;
      type_cast_778_inst_ack_1<= rack(0);
      type_cast_778_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_778_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_777_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_779,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_806_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_806_inst_req_0;
      type_cast_806_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_806_inst_req_1;
      type_cast_806_inst_ack_1<= rack(0);
      type_cast_806_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_806_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_805_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp402_807,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_822_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_822_inst_req_0;
      type_cast_822_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_822_inst_req_1;
      type_cast_822_inst_ack_1<= rack(0);
      type_cast_822_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_822_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_605,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp20_823,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_831_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_831_inst_req_0;
      type_cast_831_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_831_inst_req_1;
      type_cast_831_inst_ack_1<= rack(0);
      type_cast_831_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_831_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_630,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp22_832,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_841_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_841_inst_req_0;
      type_cast_841_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_841_inst_req_1;
      type_cast_841_inst_ack_1<= rack(0);
      type_cast_841_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_841_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_840_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp24_842,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_870_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_870_inst_req_0;
      type_cast_870_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_870_inst_req_1;
      type_cast_870_inst_ack_1<= rack(0);
      type_cast_870_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_870_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext410_1021,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_870_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_884_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_884_inst_req_0;
      type_cast_884_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_884_inst_req_1;
      type_cast_884_inst_ack_1<= rack(0);
      type_cast_884_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_884_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call89_881,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_885,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_897_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_897_inst_req_0;
      type_cast_897_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_897_inst_req_1;
      type_cast_897_inst_ack_1<= rack(0);
      type_cast_897_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_897_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call93_894,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_898,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_915_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_915_inst_req_0;
      type_cast_915_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_915_inst_req_1;
      type_cast_915_inst_ack_1<= rack(0);
      type_cast_915_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_915_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call99_912,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv101_916,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_933_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_933_inst_req_0;
      type_cast_933_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_933_inst_req_1;
      type_cast_933_inst_ack_1<= rack(0);
      type_cast_933_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_933_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call105_930,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_934,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_951_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_951_inst_req_0;
      type_cast_951_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_951_inst_req_1;
      type_cast_951_inst_ack_1<= rack(0);
      type_cast_951_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_951_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call111_948,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_952,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_969_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_969_inst_req_0;
      type_cast_969_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_969_inst_req_1;
      type_cast_969_inst_ack_1<= rack(0);
      type_cast_969_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_969_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call117_966,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv119_970,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_987_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_987_inst_req_0;
      type_cast_987_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_987_inst_req_1;
      type_cast_987_inst_ack_1<= rack(0);
      type_cast_987_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_987_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call123_984,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_988,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1192_index_1_rename
    process(R_ix_x0x_xlcssa_1191_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0x_xlcssa_1191_resized;
      ov(13 downto 0) := iv;
      R_ix_x0x_xlcssa_1191_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1192_index_1_resize
    process(ix_x0x_xlcssa_1058) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0x_xlcssa_1058;
      ov := iv(13 downto 0);
      R_ix_x0x_xlcssa_1191_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1192_root_address_inst
    process(array_obj_ref_1192_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1192_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1192_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1337_index_1_rename
    process(R_indvar395_1336_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar395_1336_resized;
      ov(13 downto 0) := iv;
      R_indvar395_1336_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1337_index_1_resize
    process(indvar395_1325) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar395_1325;
      ov := iv(13 downto 0);
      R_indvar395_1336_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1337_root_address_inst
    process(array_obj_ref_1337_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1337_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1337_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1657_index_1_rename
    process(R_ix_x1x_xlcssa_1656_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x1x_xlcssa_1656_resized;
      ov(13 downto 0) := iv;
      R_ix_x1x_xlcssa_1656_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1657_index_1_resize
    process(ix_x1x_xlcssa_1519) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x1x_xlcssa_1519;
      ov := iv(13 downto 0);
      R_ix_x1x_xlcssa_1656_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1657_root_address_inst
    process(array_obj_ref_1657_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1657_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1657_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_876_index_1_rename
    process(R_indvar409_875_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar409_875_resized;
      ov(13 downto 0) := iv;
      R_indvar409_875_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_876_index_1_resize
    process(indvar409_864) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar409_864;
      ov := iv(13 downto 0);
      R_indvar409_875_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_876_root_address_inst
    process(array_obj_ref_876_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_876_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_876_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1013_addr_0
    process(ptr_deref_1013_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1013_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1013_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1013_base_resize
    process(arrayidx_878) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_878;
      ov := iv(13 downto 0);
      ptr_deref_1013_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1013_gather_scatter
    process(add132_1011) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add132_1011;
      ov(63 downto 0) := iv;
      ptr_deref_1013_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1013_root_address_inst
    process(ptr_deref_1013_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1013_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1013_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1196_addr_0
    process(ptr_deref_1196_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1196_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1196_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1196_base_resize
    process(arrayidx143_1194) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx143_1194;
      ov := iv(13 downto 0);
      ptr_deref_1196_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1196_gather_scatter
    process(shl14x_xi_1187) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl14x_xi_1187;
      ov(63 downto 0) := iv;
      ptr_deref_1196_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1196_root_address_inst
    process(ptr_deref_1196_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1196_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1196_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1474_addr_0
    process(ptr_deref_1474_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1474_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1474_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1474_base_resize
    process(arrayidx211_1339) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx211_1339;
      ov := iv(13 downto 0);
      ptr_deref_1474_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1474_gather_scatter
    process(add207_1472) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add207_1472;
      ov(63 downto 0) := iv;
      ptr_deref_1474_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1474_root_address_inst
    process(ptr_deref_1474_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1474_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1474_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1661_addr_0
    process(ptr_deref_1661_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1661_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1661_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1661_base_resize
    process(arrayidx226_1659) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx226_1659;
      ov := iv(13 downto 0);
      ptr_deref_1661_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1661_gather_scatter
    process(shl14x_xi356_1652) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl14x_xi356_1652;
      ov(63 downto 0) := iv;
      ptr_deref_1661_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1661_root_address_inst
    process(ptr_deref_1661_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1661_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1661_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1027_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond28_1026;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1027_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1027_branch_req_0,
          ack0 => if_stmt_1027_branch_ack_0,
          ack1 => if_stmt_1027_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1078_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_1077;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1078_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1078_branch_req_0,
          ack0 => if_stmt_1078_branch_ack_0,
          ack1 => if_stmt_1078_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1153_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi_1152;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1153_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1153_branch_req_0,
          ack0 => if_stmt_1153_branch_ack_0,
          ack1 => if_stmt_1153_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1249_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp161363_1248;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1249_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1249_branch_req_0,
          ack0 => if_stmt_1249_branch_ack_0,
          ack1 => if_stmt_1249_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1488_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1487;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1488_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1488_branch_req_0,
          ack0 => if_stmt_1488_branch_ack_0,
          ack1 => if_stmt_1488_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1539_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool218_1538;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1539_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1539_branch_req_0,
          ack0 => if_stmt_1539_branch_ack_0,
          ack1 => if_stmt_1539_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1618_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi348_1617;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1618_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1618_branch_req_0,
          ack0 => if_stmt_1618_branch_ack_0,
          ack1 => if_stmt_1618_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1753_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond5_1752;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1753_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1753_branch_req_0,
          ack0 => if_stmt_1753_branch_ack_0,
          ack1 => if_stmt_1753_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_786_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp367_785;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_786_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_786_branch_req_0,
          ack0 => if_stmt_786_branch_ack_0,
          ack1 => if_stmt_786_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1118_inst
    process(nx_x022x_xi_1099) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi_1099, type_cast_1117_wire_constant, tmp_var);
      tmp_1119 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1124_inst
    process(nx_x022x_xi_1099) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi_1099, type_cast_1123_wire_constant, tmp_var);
      iNsTr_35_1125 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1583_inst
    process(nx_x022x_xi341_1564) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi341_1564, type_cast_1582_wire_constant, tmp_var);
      tmp372_1584 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1589_inst
    process(nx_x022x_xi341_1564) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi341_1564, type_cast_1588_wire_constant, tmp_var);
      iNsTr_67_1590 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1682_inst
    process(add53_705) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add53_705, type_cast_1681_wire_constant, tmp_var);
      tmp373_1683 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1020_inst
    process(indvar409_864) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar409_864, type_cast_1019_wire_constant, tmp_var);
      indvarx_xnext410_1021 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1481_inst
    process(indvar395_1325) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar395_1325, type_cast_1480_wire_constant, tmp_var);
      indvarx_xnext396_1482 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1697_inst
    process(tmp3_1692) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_1692, type_cast_1696_wire_constant, tmp_var);
      tmp4_1698 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1746_inst
    process(indvar_1710) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1710, type_cast_1745_wire_constant, tmp_var);
      indvarx_xnext_1747 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1095_inst
    process(conv2x_xi_1090) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi_1090, type_cast_1094_wire_constant, tmp_var);
      shlx_xi_1096 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1560_inst
    process(conv2x_xi338_1555) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi338_1555, type_cast_1559_wire_constant, tmp_var);
      shlx_xi339_1561 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1070_inst
    process(conv83_779) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv83_779, type_cast_1069_wire_constant, tmp_var);
      and_1071 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1175_inst
    process(Bx_xnot_1170) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(Bx_xnot_1170, type_cast_1174_wire_constant, tmp_var);
      add1216x_xi_1176 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1531_inst
    process(conv155_1242) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv155_1242, type_cast_1530_wire_constant, tmp_var);
      and217_1532 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1640_inst
    process(iNsTr_90_1635) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_90_1635, type_cast_1639_wire_constant, tmp_var);
      add1216x_xi354_1641 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1733_inst
    process(mul250_1722) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mul250_1722, type_cast_1732_wire_constant, tmp_var);
      conv251_1734 <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1053_inst
    process(type_cast_1049_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1049_wire, type_cast_1052_wire_constant, tmp_var);
      ASHR_i64_i64_1053_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1240_inst
    process(type_cast_1236_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1236_wire, type_cast_1239_wire_constant, tmp_var);
      ASHR_i64_i64_1240_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1514_inst
    process(type_cast_1510_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1510_wire, type_cast_1513_wire_constant, tmp_var);
      ASHR_i64_i64_1514_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1025_inst
    process(indvarx_xnext410_1021, umax27_861) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext410_1021, umax27_861, tmp_var);
      exitcond28_1026 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1076_inst
    process(and_1071) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and_1071, type_cast_1075_wire_constant, tmp_var);
      tobool_1077 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1486_inst
    process(indvarx_xnext396_1482, umax19_1322) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext396_1482, umax19_1322, tmp_var);
      exitcond_1487 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1537_inst
    process(and217_1532) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and217_1532, type_cast_1536_wire_constant, tmp_var);
      tobool218_1538 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1751_inst
    process(indvarx_xnext_1747, tmp4_1698) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1747, tmp4_1698, tmp_var);
      exitcond5_1752 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1260_inst
    process(conv155_1242) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv155_1242, type_cast_1259_wire_constant, tmp_var);
      tmp390_1261 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1308_inst
    process(tmp16_1303) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp16_1303, type_cast_1307_wire_constant, tmp_var);
      tmp17_1309 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1789_inst
    process(sub_1780) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1780, type_cast_1788_wire_constant, tmp_var);
      shr280_1790 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1799_inst
    process(sub_1780) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1780, type_cast_1798_wire_constant, tmp_var);
      shr286_1800 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1809_inst
    process(sub_1780) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1780, type_cast_1808_wire_constant, tmp_var);
      shr292_1810 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1819_inst
    process(sub_1780) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1780, type_cast_1818_wire_constant, tmp_var);
      shr298_1820 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1829_inst
    process(sub_1780) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1780, type_cast_1828_wire_constant, tmp_var);
      shr304_1830 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1839_inst
    process(sub_1780) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1780, type_cast_1838_wire_constant, tmp_var);
      shr310_1840 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1849_inst
    process(sub_1780) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1780, type_cast_1848_wire_constant, tmp_var);
      shr316_1850 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_812_inst
    process(tmp402_807) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp402_807, type_cast_811_wire_constant, tmp_var);
      tmp403_813 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_847_inst
    process(tmp24_842) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp24_842, type_cast_846_wire_constant, tmp_var);
      tmp25_848 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1687_inst
    process(add73_755, add23_630) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_755, add23_630, tmp_var);
      tmp377_1688 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_767_inst
    process(conv79_759, add_580) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv79_759, add_580, tmp_var);
      mul_768 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_772_inst
    process(mul_768, conv81_763) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_768, conv81_763, tmp_var);
      mul82_773 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_796_inst
    process(add_580, conv79_759) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_580, conv79_759, tmp_var);
      tmp399_797 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_801_inst
    process(tmp399_797, conv81_763) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp399_797, conv81_763, tmp_var);
      tmp401_802 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_827_inst
    process(add_580, tmp20_823) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_580, tmp20_823, tmp_var);
      tmp21_828 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_836_inst
    process(tmp21_828, tmp22_832) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp21_828, tmp22_832, tmp_var);
      tmp23_837 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1216_inst
    process(conv153_1212, conv145_1204) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv153_1212, conv145_1204, tmp_var);
      mul148_1217 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1221_inst
    process(mul148_1217, add63_730) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul148_1217, add63_730, tmp_var);
      mul151_1222 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1226_inst
    process(mul151_1222, conv147_1208) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul151_1222, conv147_1208, tmp_var);
      mul154_1227 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1275_inst
    process(add63_730, tmp9_1271) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add63_730, tmp9_1271, tmp_var);
      tmp10_1276 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1284_inst
    process(tmp10_1276, tmp11_1280) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp10_1276, tmp11_1280, tmp_var);
      tmp12_1285 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1293_inst
    process(tmp12_1285, tmp13_1289) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp12_1285, tmp13_1289, tmp_var);
      tmp14_1294 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1706_inst
    process(add63_730, tmp6_1702) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(add63_730, tmp6_1702, tmp_var);
      tmp7_1707 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1721_inst
    process(tmp7_1707, indvar_1710) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp7_1707, indvar_1710, tmp_var);
      mul250_1722 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_604_inst
    process(shl10_593, conv12_600) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl10_593, conv12_600, tmp_var);
      add13_605 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_629_inst
    process(shl20_618, conv22_625) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl20_618, conv22_625, tmp_var);
      add23_630 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_654_inst
    process(shl30_643, conv32_650) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl30_643, conv32_650, tmp_var);
      add33_655 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_679_inst
    process(shl40_668, conv42_675) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl40_668, conv42_675, tmp_var);
      add43_680 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_704_inst
    process(shl50_693, conv52_700) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl50_693, conv52_700, tmp_var);
      add53_705 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_754_inst
    process(shl70_743, conv72_750) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl70_743, conv72_750, tmp_var);
      add73_755 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_579_inst
    process(shl_568, conv3_575) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_568, conv3_575, tmp_var);
      add_580 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1010_inst
    process(shl128_999, conv131_1006) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl128_999, conv131_1006, tmp_var);
      add132_1011 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1136_inst
    process(conv5x_xi_1132, elementx_x021x_xi_1106) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi_1132, elementx_x021x_xi_1106, tmp_var);
      addx_xi_1137 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1363_inst
    process(shl167_1352, conv170_1359) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl167_1352, conv170_1359, tmp_var);
      add171_1364 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1381_inst
    process(shl173_1370, conv176_1377) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl173_1370, conv176_1377, tmp_var);
      add177_1382 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1399_inst
    process(shl179_1388, conv182_1395) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl179_1388, conv182_1395, tmp_var);
      add183_1400 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1417_inst
    process(shl185_1406, conv188_1413) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl185_1406, conv188_1413, tmp_var);
      add189_1418 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1435_inst
    process(shl191_1424, conv194_1431) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl191_1424, conv194_1431, tmp_var);
      add195_1436 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1453_inst
    process(shl197_1442, conv200_1449) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl197_1442, conv200_1449, tmp_var);
      add201_1454 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1471_inst
    process(shl203_1460, conv206_1467) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl203_1460, conv206_1467, tmp_var);
      add207_1472 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1601_inst
    process(conv5x_xi344_1597, elementx_x021x_xi342_1571) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi344_1597, elementx_x021x_xi342_1571, tmp_var);
      addx_xi345_1602 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_729_inst
    process(shl60_718, conv62_725) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl60_718, conv62_725, tmp_var);
      add63_730 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_902_inst
    process(shl92_891, conv95_898) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl92_891, conv95_898, tmp_var);
      add96_903 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_920_inst
    process(shl98_909, conv101_916) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl98_909, conv101_916, tmp_var);
      add102_921 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_938_inst
    process(shl104_927, conv107_934) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl104_927, conv107_934, tmp_var);
      add108_939 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_956_inst
    process(shl110_945, conv113_952) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl110_945, conv113_952, tmp_var);
      add114_957 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_974_inst
    process(shl116_963, conv119_970) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl116_963, conv119_970, tmp_var);
      add120_975 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_992_inst
    process(shl122_981, conv125_988) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl122_981, conv125_988, tmp_var);
      add126_993 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_592_inst
    process(conv9_587) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv9_587, type_cast_591_wire_constant, tmp_var);
      shl10_593 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_617_inst
    process(conv19_612) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_612, type_cast_616_wire_constant, tmp_var);
      shl20_618 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_642_inst
    process(conv29_637) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv29_637, type_cast_641_wire_constant, tmp_var);
      shl30_643 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_667_inst
    process(conv39_662) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv39_662, type_cast_666_wire_constant, tmp_var);
      shl40_668 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_692_inst
    process(conv49_687) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_687, type_cast_691_wire_constant, tmp_var);
      shl50_693 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_742_inst
    process(conv69_737) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv69_737, type_cast_741_wire_constant, tmp_var);
      shl70_743 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1089_inst
    process(mul82_773) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul82_773, type_cast_1088_wire_constant, tmp_var);
      conv2x_xi_1090 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_567_inst
    process(conv1_562) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_562, type_cast_566_wire_constant, tmp_var);
      shl_568 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1045_inst
    process(umax405_1040) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax405_1040, type_cast_1044_wire_constant, tmp_var);
      tmp406_1046 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1142_inst
    process(addx_xi_1137) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi_1137, type_cast_1141_wire_constant, tmp_var);
      shl8x_xi_1143 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1169_inst
    process(conv83_779) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv83_779, type_cast_1168_wire_constant, tmp_var);
      Bx_xnot_1170 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1186_inst
    process(shl8x_xix_xlcssa_1160, sh_promx_xi_1182) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl8x_xix_xlcssa_1160, sh_promx_xi_1182, tmp_var);
      shl14x_xi_1187 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1232_inst
    process(mul154_1227) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1227, type_cast_1231_wire_constant, tmp_var);
      sext_1233 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1351_inst
    process(conv165_1346) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv165_1346, type_cast_1350_wire_constant, tmp_var);
      shl167_1352 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1369_inst
    process(add171_1364) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add171_1364, type_cast_1368_wire_constant, tmp_var);
      shl173_1370 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1387_inst
    process(add177_1382) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add177_1382, type_cast_1386_wire_constant, tmp_var);
      shl179_1388 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1405_inst
    process(add183_1400) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add183_1400, type_cast_1404_wire_constant, tmp_var);
      shl185_1406 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1423_inst
    process(add189_1418) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add189_1418, type_cast_1422_wire_constant, tmp_var);
      shl191_1424 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1441_inst
    process(add195_1436) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add195_1436, type_cast_1440_wire_constant, tmp_var);
      shl197_1442 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1459_inst
    process(add201_1454) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add201_1454, type_cast_1458_wire_constant, tmp_var);
      shl203_1460 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1506_inst
    process(umax_1501) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax_1501, type_cast_1505_wire_constant, tmp_var);
      tmp392_1507 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1550_inst
    process(mul154_1227) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1227, type_cast_1549_wire_constant, tmp_var);
      iNsTr_55_1551 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1607_inst
    process(addx_xi345_1602) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi345_1602, type_cast_1606_wire_constant, tmp_var);
      shl8x_xi346_1608 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1634_inst
    process(mul154_1227) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1227, type_cast_1633_wire_constant, tmp_var);
      iNsTr_90_1635 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1651_inst
    process(shl8x_xi346x_xlcssa_1625, sh_promx_xi355_1647) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl8x_xi346x_xlcssa_1625, sh_promx_xi355_1647, tmp_var);
      shl14x_xi356_1652 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_717_inst
    process(conv59_712) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv59_712, type_cast_716_wire_constant, tmp_var);
      shl60_718 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_890_inst
    process(conv90_885) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv90_885, type_cast_889_wire_constant, tmp_var);
      shl92_891 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_908_inst
    process(add96_903) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add96_903, type_cast_907_wire_constant, tmp_var);
      shl98_909 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_926_inst
    process(add102_921) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add102_921, type_cast_925_wire_constant, tmp_var);
      shl104_927 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_944_inst
    process(add108_939) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add108_939, type_cast_943_wire_constant, tmp_var);
      shl110_945 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_962_inst
    process(add114_957) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add114_957, type_cast_961_wire_constant, tmp_var);
      shl116_963 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_980_inst
    process(add120_975) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add120_975, type_cast_979_wire_constant, tmp_var);
      shl122_981 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_998_inst
    process(add126_993) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add126_993, type_cast_997_wire_constant, tmp_var);
      shl128_999 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1779_inst
    process(conv270_1775, conv230_1764) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv270_1775, conv230_1764, tmp_var);
      sub_1780 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_784_inst
    process(mul82_773) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul82_773, type_cast_783_wire_constant, tmp_var);
      cmp367_785 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1247_inst
    process(conv155_1242) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv155_1242, type_cast_1246_wire_constant, tmp_var);
      cmp161363_1248 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1266_inst
    process(tmp390_1261) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp390_1261, type_cast_1265_wire_constant, tmp_var);
      tmp391_1267 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1314_inst
    process(tmp17_1309) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp17_1309, type_cast_1313_wire_constant, tmp_var);
      tmp18_1315 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_818_inst
    process(tmp403_813) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp403_813, type_cast_817_wire_constant, tmp_var);
      tmp404_819 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_853_inst
    process(tmp25_848) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp25_848, type_cast_852_wire_constant, tmp_var);
      tmp26_854 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1151_inst
    process(convx_xi_1147, shlx_xi_1096) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi_1147, shlx_xi_1096, tmp_var);
      cmpx_xi_1152 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1616_inst
    process(convx_xi347_1612, shlx_xi339_1561) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi347_1612, shlx_xi339_1561, tmp_var);
      cmpx_xi348_1617 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_1181_inst
    process(add1216x_xi_1176) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1216x_xi_1176, type_cast_1180_wire_constant, tmp_var);
      sh_promx_xi_1182 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_1646_inst
    process(add1216x_xi354_1641) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1216x_xi354_1641, type_cast_1645_wire_constant, tmp_var);
      sh_promx_xi355_1647 <= tmp_var; --
    end process;
    -- shared split operator group (118) : array_obj_ref_1192_index_offset 
    ApIntAdd_group_118: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0x_xlcssa_1191_scaled;
      array_obj_ref_1192_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1192_index_offset_req_0;
      array_obj_ref_1192_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1192_index_offset_req_1;
      array_obj_ref_1192_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_118_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_118_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_118",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 118
    -- shared split operator group (119) : array_obj_ref_1337_index_offset 
    ApIntAdd_group_119: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar395_1336_scaled;
      array_obj_ref_1337_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1337_index_offset_req_0;
      array_obj_ref_1337_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1337_index_offset_req_1;
      array_obj_ref_1337_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_119_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_119_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_119",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 119
    -- shared split operator group (120) : array_obj_ref_1657_index_offset 
    ApIntAdd_group_120: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x1x_xlcssa_1656_scaled;
      array_obj_ref_1657_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1657_index_offset_req_0;
      array_obj_ref_1657_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1657_index_offset_req_1;
      array_obj_ref_1657_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_120_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_120_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_120",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 120
    -- shared split operator group (121) : array_obj_ref_876_index_offset 
    ApIntAdd_group_121: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar409_875_scaled;
      array_obj_ref_876_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_876_index_offset_req_0;
      array_obj_ref_876_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_876_index_offset_req_1;
      array_obj_ref_876_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_121_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_121_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_121",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 121
    -- unary operator type_cast_1301_inst
    process(tmp15_1298) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp15_1298, tmp_var);
      type_cast_1301_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1762_inst
    process(call229_1668) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call229_1668, tmp_var);
      type_cast_1762_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1773_inst
    process(call269_1770) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call269_1770, tmp_var);
      type_cast_1773_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_777_inst
    process(mul82_773) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", mul82_773, tmp_var);
      type_cast_777_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_805_inst
    process(tmp401_802) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp401_802, tmp_var);
      type_cast_805_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_840_inst
    process(tmp23_837) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp23_837, tmp_var);
      type_cast_840_wire <= tmp_var; -- 
    end process;
    -- shared store operator group (0) : ptr_deref_1013_store_0 ptr_deref_1196_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1013_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1196_store_0_req_0;
      ptr_deref_1013_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1196_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1013_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1196_store_0_req_1;
      ptr_deref_1013_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1196_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1013_word_address_0 & ptr_deref_1196_word_address_0;
      data_in <= ptr_deref_1013_data_0 & ptr_deref_1196_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1474_store_0 ptr_deref_1661_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1474_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1661_store_0_req_0;
      ptr_deref_1474_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1661_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1474_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1661_store_0_req_1;
      ptr_deref_1474_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1661_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1474_word_address_0 & ptr_deref_1661_word_address_0;
      data_in <= ptr_deref_1474_data_0 & ptr_deref_1661_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : RPIPE_input_done_pipe_1766_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_done_pipe_1766_inst_req_0;
      RPIPE_input_done_pipe_1766_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_done_pipe_1766_inst_req_1;
      RPIPE_input_done_pipe_1766_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call267_1767 <= data_out(7 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_maxpool_input_pipe_947_inst RPIPE_maxpool_input_pipe_1341_inst RPIPE_maxpool_input_pipe_965_inst RPIPE_maxpool_input_pipe_983_inst RPIPE_maxpool_input_pipe_1001_inst RPIPE_maxpool_input_pipe_1354_inst RPIPE_maxpool_input_pipe_1127_inst RPIPE_maxpool_input_pipe_1408_inst RPIPE_maxpool_input_pipe_1444_inst RPIPE_maxpool_input_pipe_1390_inst RPIPE_maxpool_input_pipe_1462_inst RPIPE_maxpool_input_pipe_1372_inst RPIPE_maxpool_input_pipe_929_inst RPIPE_maxpool_input_pipe_893_inst RPIPE_maxpool_input_pipe_1426_inst RPIPE_maxpool_input_pipe_911_inst RPIPE_maxpool_input_pipe_557_inst RPIPE_maxpool_input_pipe_570_inst RPIPE_maxpool_input_pipe_582_inst RPIPE_maxpool_input_pipe_595_inst RPIPE_maxpool_input_pipe_607_inst RPIPE_maxpool_input_pipe_620_inst RPIPE_maxpool_input_pipe_632_inst RPIPE_maxpool_input_pipe_645_inst RPIPE_maxpool_input_pipe_657_inst RPIPE_maxpool_input_pipe_670_inst RPIPE_maxpool_input_pipe_682_inst RPIPE_maxpool_input_pipe_695_inst RPIPE_maxpool_input_pipe_707_inst RPIPE_maxpool_input_pipe_720_inst RPIPE_maxpool_input_pipe_732_inst RPIPE_maxpool_input_pipe_745_inst RPIPE_maxpool_input_pipe_880_inst RPIPE_maxpool_input_pipe_1592_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(271 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 33 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 33 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 33 downto 0);
      signal guard_vector : std_logic_vector( 33 downto 0);
      constant outBUFs : IntegerArray(33 downto 0) := (33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(33 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false);
      constant guardBuffering: IntegerArray(33 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2);
      -- 
    begin -- 
      reqL_unguarded(33) <= RPIPE_maxpool_input_pipe_947_inst_req_0;
      reqL_unguarded(32) <= RPIPE_maxpool_input_pipe_1341_inst_req_0;
      reqL_unguarded(31) <= RPIPE_maxpool_input_pipe_965_inst_req_0;
      reqL_unguarded(30) <= RPIPE_maxpool_input_pipe_983_inst_req_0;
      reqL_unguarded(29) <= RPIPE_maxpool_input_pipe_1001_inst_req_0;
      reqL_unguarded(28) <= RPIPE_maxpool_input_pipe_1354_inst_req_0;
      reqL_unguarded(27) <= RPIPE_maxpool_input_pipe_1127_inst_req_0;
      reqL_unguarded(26) <= RPIPE_maxpool_input_pipe_1408_inst_req_0;
      reqL_unguarded(25) <= RPIPE_maxpool_input_pipe_1444_inst_req_0;
      reqL_unguarded(24) <= RPIPE_maxpool_input_pipe_1390_inst_req_0;
      reqL_unguarded(23) <= RPIPE_maxpool_input_pipe_1462_inst_req_0;
      reqL_unguarded(22) <= RPIPE_maxpool_input_pipe_1372_inst_req_0;
      reqL_unguarded(21) <= RPIPE_maxpool_input_pipe_929_inst_req_0;
      reqL_unguarded(20) <= RPIPE_maxpool_input_pipe_893_inst_req_0;
      reqL_unguarded(19) <= RPIPE_maxpool_input_pipe_1426_inst_req_0;
      reqL_unguarded(18) <= RPIPE_maxpool_input_pipe_911_inst_req_0;
      reqL_unguarded(17) <= RPIPE_maxpool_input_pipe_557_inst_req_0;
      reqL_unguarded(16) <= RPIPE_maxpool_input_pipe_570_inst_req_0;
      reqL_unguarded(15) <= RPIPE_maxpool_input_pipe_582_inst_req_0;
      reqL_unguarded(14) <= RPIPE_maxpool_input_pipe_595_inst_req_0;
      reqL_unguarded(13) <= RPIPE_maxpool_input_pipe_607_inst_req_0;
      reqL_unguarded(12) <= RPIPE_maxpool_input_pipe_620_inst_req_0;
      reqL_unguarded(11) <= RPIPE_maxpool_input_pipe_632_inst_req_0;
      reqL_unguarded(10) <= RPIPE_maxpool_input_pipe_645_inst_req_0;
      reqL_unguarded(9) <= RPIPE_maxpool_input_pipe_657_inst_req_0;
      reqL_unguarded(8) <= RPIPE_maxpool_input_pipe_670_inst_req_0;
      reqL_unguarded(7) <= RPIPE_maxpool_input_pipe_682_inst_req_0;
      reqL_unguarded(6) <= RPIPE_maxpool_input_pipe_695_inst_req_0;
      reqL_unguarded(5) <= RPIPE_maxpool_input_pipe_707_inst_req_0;
      reqL_unguarded(4) <= RPIPE_maxpool_input_pipe_720_inst_req_0;
      reqL_unguarded(3) <= RPIPE_maxpool_input_pipe_732_inst_req_0;
      reqL_unguarded(2) <= RPIPE_maxpool_input_pipe_745_inst_req_0;
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_880_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_1592_inst_req_0;
      RPIPE_maxpool_input_pipe_947_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_maxpool_input_pipe_1341_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_maxpool_input_pipe_965_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_maxpool_input_pipe_983_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_maxpool_input_pipe_1001_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_maxpool_input_pipe_1354_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_maxpool_input_pipe_1127_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_maxpool_input_pipe_1408_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_maxpool_input_pipe_1444_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_maxpool_input_pipe_1390_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_maxpool_input_pipe_1462_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_maxpool_input_pipe_1372_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_maxpool_input_pipe_929_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_maxpool_input_pipe_893_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_maxpool_input_pipe_1426_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_maxpool_input_pipe_911_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_maxpool_input_pipe_557_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_maxpool_input_pipe_570_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_maxpool_input_pipe_582_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_maxpool_input_pipe_595_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_maxpool_input_pipe_607_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_maxpool_input_pipe_620_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_maxpool_input_pipe_632_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_maxpool_input_pipe_645_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_maxpool_input_pipe_657_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_maxpool_input_pipe_670_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_maxpool_input_pipe_682_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_maxpool_input_pipe_695_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_maxpool_input_pipe_707_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_maxpool_input_pipe_720_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_maxpool_input_pipe_732_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_maxpool_input_pipe_745_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_maxpool_input_pipe_880_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_1592_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(33) <= RPIPE_maxpool_input_pipe_947_inst_req_1;
      reqR_unguarded(32) <= RPIPE_maxpool_input_pipe_1341_inst_req_1;
      reqR_unguarded(31) <= RPIPE_maxpool_input_pipe_965_inst_req_1;
      reqR_unguarded(30) <= RPIPE_maxpool_input_pipe_983_inst_req_1;
      reqR_unguarded(29) <= RPIPE_maxpool_input_pipe_1001_inst_req_1;
      reqR_unguarded(28) <= RPIPE_maxpool_input_pipe_1354_inst_req_1;
      reqR_unguarded(27) <= RPIPE_maxpool_input_pipe_1127_inst_req_1;
      reqR_unguarded(26) <= RPIPE_maxpool_input_pipe_1408_inst_req_1;
      reqR_unguarded(25) <= RPIPE_maxpool_input_pipe_1444_inst_req_1;
      reqR_unguarded(24) <= RPIPE_maxpool_input_pipe_1390_inst_req_1;
      reqR_unguarded(23) <= RPIPE_maxpool_input_pipe_1462_inst_req_1;
      reqR_unguarded(22) <= RPIPE_maxpool_input_pipe_1372_inst_req_1;
      reqR_unguarded(21) <= RPIPE_maxpool_input_pipe_929_inst_req_1;
      reqR_unguarded(20) <= RPIPE_maxpool_input_pipe_893_inst_req_1;
      reqR_unguarded(19) <= RPIPE_maxpool_input_pipe_1426_inst_req_1;
      reqR_unguarded(18) <= RPIPE_maxpool_input_pipe_911_inst_req_1;
      reqR_unguarded(17) <= RPIPE_maxpool_input_pipe_557_inst_req_1;
      reqR_unguarded(16) <= RPIPE_maxpool_input_pipe_570_inst_req_1;
      reqR_unguarded(15) <= RPIPE_maxpool_input_pipe_582_inst_req_1;
      reqR_unguarded(14) <= RPIPE_maxpool_input_pipe_595_inst_req_1;
      reqR_unguarded(13) <= RPIPE_maxpool_input_pipe_607_inst_req_1;
      reqR_unguarded(12) <= RPIPE_maxpool_input_pipe_620_inst_req_1;
      reqR_unguarded(11) <= RPIPE_maxpool_input_pipe_632_inst_req_1;
      reqR_unguarded(10) <= RPIPE_maxpool_input_pipe_645_inst_req_1;
      reqR_unguarded(9) <= RPIPE_maxpool_input_pipe_657_inst_req_1;
      reqR_unguarded(8) <= RPIPE_maxpool_input_pipe_670_inst_req_1;
      reqR_unguarded(7) <= RPIPE_maxpool_input_pipe_682_inst_req_1;
      reqR_unguarded(6) <= RPIPE_maxpool_input_pipe_695_inst_req_1;
      reqR_unguarded(5) <= RPIPE_maxpool_input_pipe_707_inst_req_1;
      reqR_unguarded(4) <= RPIPE_maxpool_input_pipe_720_inst_req_1;
      reqR_unguarded(3) <= RPIPE_maxpool_input_pipe_732_inst_req_1;
      reqR_unguarded(2) <= RPIPE_maxpool_input_pipe_745_inst_req_1;
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_880_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_1592_inst_req_1;
      RPIPE_maxpool_input_pipe_947_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_maxpool_input_pipe_1341_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_maxpool_input_pipe_965_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_maxpool_input_pipe_983_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_maxpool_input_pipe_1001_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_maxpool_input_pipe_1354_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_maxpool_input_pipe_1127_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_maxpool_input_pipe_1408_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_maxpool_input_pipe_1444_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_maxpool_input_pipe_1390_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_maxpool_input_pipe_1462_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_maxpool_input_pipe_1372_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_maxpool_input_pipe_929_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_maxpool_input_pipe_893_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_maxpool_input_pipe_1426_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_maxpool_input_pipe_911_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_maxpool_input_pipe_557_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_maxpool_input_pipe_570_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_maxpool_input_pipe_582_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_maxpool_input_pipe_595_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_maxpool_input_pipe_607_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_maxpool_input_pipe_620_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_maxpool_input_pipe_632_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_maxpool_input_pipe_645_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_maxpool_input_pipe_657_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_maxpool_input_pipe_670_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_maxpool_input_pipe_682_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_maxpool_input_pipe_695_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_maxpool_input_pipe_707_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_maxpool_input_pipe_720_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_maxpool_input_pipe_732_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_maxpool_input_pipe_745_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_maxpool_input_pipe_880_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_1592_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      call111_948 <= data_out(271 downto 264);
      call164_1342 <= data_out(263 downto 256);
      call117_966 <= data_out(255 downto 248);
      call123_984 <= data_out(247 downto 240);
      call129_1002 <= data_out(239 downto 232);
      call168_1355 <= data_out(231 downto 224);
      callx_xi_1128 <= data_out(223 downto 216);
      call186_1409 <= data_out(215 downto 208);
      call198_1445 <= data_out(207 downto 200);
      call180_1391 <= data_out(199 downto 192);
      call204_1463 <= data_out(191 downto 184);
      call174_1373 <= data_out(183 downto 176);
      call105_930 <= data_out(175 downto 168);
      call93_894 <= data_out(167 downto 160);
      call192_1427 <= data_out(159 downto 152);
      call99_912 <= data_out(151 downto 144);
      call_558 <= data_out(143 downto 136);
      call2_571 <= data_out(135 downto 128);
      call6_583 <= data_out(127 downto 120);
      call11_596 <= data_out(119 downto 112);
      call16_608 <= data_out(111 downto 104);
      call21_621 <= data_out(103 downto 96);
      call26_633 <= data_out(95 downto 88);
      call31_646 <= data_out(87 downto 80);
      call36_658 <= data_out(79 downto 72);
      call41_671 <= data_out(71 downto 64);
      call46_683 <= data_out(63 downto 56);
      call51_696 <= data_out(55 downto 48);
      call56_708 <= data_out(47 downto 40);
      call61_721 <= data_out(39 downto 32);
      call66_733 <= data_out(31 downto 24);
      call71_746 <= data_out(23 downto 16);
      call89_881 <= data_out(15 downto 8);
      callx_xi343_1593 <= data_out(7 downto 0);
      maxpool_input_pipe_read_1_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_1_gI", nreqs => 34, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_1: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_1", data_width => 8,  num_reqs => 34,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_1670_inst WPIPE_maxpool_output_pipe_1674_inst WPIPE_maxpool_output_pipe_1855_inst WPIPE_maxpool_output_pipe_1858_inst WPIPE_maxpool_output_pipe_1861_inst WPIPE_maxpool_output_pipe_1864_inst WPIPE_maxpool_output_pipe_1867_inst WPIPE_maxpool_output_pipe_1870_inst WPIPE_maxpool_output_pipe_1873_inst WPIPE_maxpool_output_pipe_1876_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal sample_req, sample_ack : BooleanArray( 9 downto 0);
      signal update_req, update_ack : BooleanArray( 9 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 9 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 9 downto 0);
      signal guard_vector : std_logic_vector( 9 downto 0);
      constant inBUFs : IntegerArray(9 downto 0) := (9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(9 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false);
      constant guardBuffering: IntegerArray(9 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2);
      -- 
    begin -- 
      sample_req_unguarded(9) <= WPIPE_maxpool_output_pipe_1670_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_maxpool_output_pipe_1674_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_1855_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_1858_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1861_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_1864_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1867_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1870_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1873_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1876_inst_req_0;
      WPIPE_maxpool_output_pipe_1670_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_maxpool_output_pipe_1674_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_maxpool_output_pipe_1855_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_1858_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1861_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_1864_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1867_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1870_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1873_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1876_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(9) <= WPIPE_maxpool_output_pipe_1670_inst_req_1;
      update_req_unguarded(8) <= WPIPE_maxpool_output_pipe_1674_inst_req_1;
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_1855_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_1858_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1861_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_1864_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1867_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1870_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1873_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1876_inst_req_1;
      WPIPE_maxpool_output_pipe_1670_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_maxpool_output_pipe_1674_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_maxpool_output_pipe_1855_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_1858_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1861_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_1864_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1867_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1870_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1873_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1876_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      data_in <= type_cast_1672_wire_constant & type_cast_1676_wire_constant & conv319_1854 & conv313_1844 & conv307_1834 & conv301_1824 & conv295_1814 & conv289_1804 & conv283_1794 & conv277_1784;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 10, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 10, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_num_out_pipe_1723_inst WPIPE_num_out_pipe_1726_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_num_out_pipe_1723_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_num_out_pipe_1726_inst_req_0;
      WPIPE_num_out_pipe_1723_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_num_out_pipe_1726_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_num_out_pipe_1723_inst_req_1;
      update_req_unguarded(0) <= WPIPE_num_out_pipe_1726_inst_req_1;
      WPIPE_num_out_pipe_1723_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_num_out_pipe_1726_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      data_in <= add33_655 & add43_680;
      num_out_pipe_write_1_gI: SplitGuardInterface generic map(name => "num_out_pipe_write_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "num_out_pipe", data_width => 16, num_reqs => 2, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => num_out_pipe_pipe_write_req(0),
          oack => num_out_pipe_pipe_write_ack(0),
          odata => num_out_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_1668_call call_stmt_1770_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1668_call_req_0;
      reqL_unguarded(0) <= call_stmt_1770_call_req_0;
      call_stmt_1668_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1770_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1668_call_req_1;
      reqR_unguarded(0) <= call_stmt_1770_call_req_1;
      call_stmt_1668_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1770_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call229_1668 <= data_out(127 downto 64);
      call269_1770 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1737_call 
    loadKernelChannel_call_group_1: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1737_call_req_0;
      call_stmt_1737_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1737_call_req_1;
      call_stmt_1737_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadKernelChannel_call_group_1_gI: SplitGuardInterface generic map(name => "loadKernelChannel_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= conv251_1734 & add23_630;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 80,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadKernelChannel_call_reqs(0),
          ackR => loadKernelChannel_call_acks(0),
          dataR => loadKernelChannel_call_data(79 downto 0),
          tagR => loadKernelChannel_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => loadKernelChannel_return_acks(0), -- cross-over
          ackL => loadKernelChannel_return_reqs(0), -- cross-over
          tagL => loadKernelChannel_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1741_call 
    access_T_call_group_2: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1741_call_req_0;
      call_stmt_1741_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1741_call_req_1;
      call_stmt_1741_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      access_T_call_group_2_gI: SplitGuardInterface generic map(name => "access_T_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= add33_655 & add23_630 & add13_605;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 48,
        owidth => 48,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => access_T_call_reqs(0),
          ackR => access_T_call_acks(0),
          dataR => access_T_call_data(47 downto 0),
          tagR => access_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => access_T_return_acks(0), -- cross-over
          ackL => access_T_return_reqs(0), -- cross-over
          tagL => access_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end convolution3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolve is -- 
  generic (tag_length : integer); 
  port ( -- 
    input_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe3_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    kernel_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
    kernel_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_read_data : in   std_logic_vector(15 downto 0);
    kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolve;
architecture convolve_arch of convolve is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolve_CP_4643_start: Boolean;
  signal convolve_CP_4643_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal phi_stmt_1926_req_1 : boolean;
  signal n_col_2230_1925_buf_ack_0 : boolean;
  signal n_row_2238_1920_buf_ack_1 : boolean;
  signal phi_stmt_1910_req_0 : boolean;
  signal n_row_2238_1920_buf_req_1 : boolean;
  signal phi_stmt_1926_req_0 : boolean;
  signal phi_stmt_1910_req_1 : boolean;
  signal do_while_stmt_1908_branch_req_0 : boolean;
  signal slice_2254_inst_req_0 : boolean;
  signal slice_2254_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_2198_inst_req_0 : boolean;
  signal slice_2254_inst_ack_1 : boolean;
  signal W_read_k_2017_delayed_1_0_2082_inst_ack_1 : boolean;
  signal W_read_k_2017_delayed_1_0_2082_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_2198_inst_ack_0 : boolean;
  signal slice_2254_inst_ack_0 : boolean;
  signal n_col_2230_1925_buf_req_1 : boolean;
  signal phi_stmt_1916_req_1 : boolean;
  signal n_chl_2208_1936_buf_ack_0 : boolean;
  signal W_store_kernel_2113_delayed_1_0_2194_inst_ack_1 : boolean;
  signal nacc_2247_1915_buf_req_0 : boolean;
  signal n_col_2230_1925_buf_ack_1 : boolean;
  signal nacc_2247_1915_buf_ack_0 : boolean;
  signal phi_stmt_1910_ack_0 : boolean;
  signal n_chl_2208_1936_buf_req_0 : boolean;
  signal n_num_2219_1931_buf_req_0 : boolean;
  signal phi_stmt_1926_ack_0 : boolean;
  signal phi_stmt_1916_req_0 : boolean;
  signal phi_stmt_1921_req_1 : boolean;
  signal n_num_2219_1931_buf_req_1 : boolean;
  signal phi_stmt_1932_ack_0 : boolean;
  signal W_acc_2059_delayed_1_0_2130_inst_req_1 : boolean;
  signal n_col_2230_1925_buf_req_0 : boolean;
  signal W_store_kernel_2113_delayed_1_0_2194_inst_req_0 : boolean;
  signal n_num_2219_1931_buf_ack_0 : boolean;
  signal phi_stmt_1921_req_0 : boolean;
  signal W_store_kernel_2105_delayed_1_0_2180_inst_ack_0 : boolean;
  signal W_acc_2059_delayed_1_0_2130_inst_ack_1 : boolean;
  signal n_num_2219_1931_buf_ack_1 : boolean;
  signal nacc_2247_1915_buf_req_1 : boolean;
  signal phi_stmt_1932_req_1 : boolean;
  signal W_store_kernel_2113_delayed_1_0_2194_inst_req_1 : boolean;
  signal nacc_2247_1915_buf_ack_1 : boolean;
  signal phi_stmt_1916_ack_0 : boolean;
  signal phi_stmt_1921_ack_0 : boolean;
  signal n_chl_2208_1936_buf_req_1 : boolean;
  signal n_chl_2208_1936_buf_ack_1 : boolean;
  signal W_num_done_2174_delayed_2_0_2264_inst_ack_1 : boolean;
  signal W_store_kernel_2113_delayed_1_0_2194_inst_ack_0 : boolean;
  signal n_row_2238_1920_buf_req_0 : boolean;
  signal phi_stmt_1932_req_0 : boolean;
  signal n_row_2238_1920_buf_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2268_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2268_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2268_inst_ack_1 : boolean;
  signal W_read_k_2017_delayed_1_0_2082_inst_req_0 : boolean;
  signal W_store_kernel_2105_delayed_1_0_2180_inst_req_1 : boolean;
  signal type_cast_2270_inst_ack_0 : boolean;
  signal W_store_kernel_2105_delayed_1_0_2180_inst_ack_1 : boolean;
  signal W_read_k_2017_delayed_1_0_2082_inst_ack_0 : boolean;
  signal type_cast_2270_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_2198_inst_req_1 : boolean;
  signal W_store_kernel_2105_delayed_1_0_2180_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_2268_inst_req_0 : boolean;
  signal W_num_done_2174_delayed_2_0_2264_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_1894_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_1894_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_1894_inst_req_1 : boolean;
  signal RPIPE_num_out_pipe_1894_inst_ack_1 : boolean;
  signal SUB_u16_u16_1896_inst_req_0 : boolean;
  signal SUB_u16_u16_1896_inst_ack_0 : boolean;
  signal SUB_u16_u16_1896_inst_req_1 : boolean;
  signal SUB_u16_u16_1896_inst_ack_1 : boolean;
  signal RPIPE_num_out_pipe_1899_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_1899_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_1899_inst_req_1 : boolean;
  signal RPIPE_num_out_pipe_1899_inst_ack_1 : boolean;
  signal SUB_u16_u16_1901_inst_req_0 : boolean;
  signal SUB_u16_u16_1901_inst_ack_0 : boolean;
  signal SUB_u16_u16_1901_inst_req_1 : boolean;
  signal SUB_u16_u16_1901_inst_ack_1 : boolean;
  signal RPIPE_size_pipe_1904_inst_req_0 : boolean;
  signal RPIPE_size_pipe_1904_inst_ack_0 : boolean;
  signal RPIPE_size_pipe_1904_inst_req_1 : boolean;
  signal RPIPE_size_pipe_1904_inst_ack_1 : boolean;
  signal SUB_u16_u16_1906_inst_req_0 : boolean;
  signal SUB_u16_u16_1906_inst_ack_0 : boolean;
  signal SUB_u16_u16_1906_inst_req_1 : boolean;
  signal SUB_u16_u16_1906_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_2184_inst_req_0 : boolean;
  signal RPIPE_input_pipe1_1949_inst_req_0 : boolean;
  signal RPIPE_input_pipe1_1949_inst_ack_0 : boolean;
  signal W_acc_2059_delayed_1_0_2130_inst_ack_0 : boolean;
  signal RPIPE_input_pipe1_1949_inst_req_1 : boolean;
  signal RPIPE_input_pipe1_1949_inst_ack_1 : boolean;
  signal W_num_done_2174_delayed_2_0_2264_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2260_inst_ack_0 : boolean;
  signal RPIPE_input_pipe2_1953_inst_req_0 : boolean;
  signal RPIPE_input_pipe2_1953_inst_ack_0 : boolean;
  signal W_acc_2059_delayed_1_0_2130_inst_req_0 : boolean;
  signal RPIPE_input_pipe2_1953_inst_req_1 : boolean;
  signal RPIPE_input_pipe2_1953_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_2191_inst_ack_1 : boolean;
  signal RPIPE_input_pipe3_1957_inst_req_0 : boolean;
  signal slice_2250_inst_ack_1 : boolean;
  signal RPIPE_input_pipe3_1957_inst_ack_0 : boolean;
  signal RPIPE_input_pipe3_1957_inst_req_1 : boolean;
  signal slice_2250_inst_req_1 : boolean;
  signal RPIPE_input_pipe3_1957_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_2191_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_2191_inst_ack_0 : boolean;
  signal W_read_k_2011_delayed_1_0_2073_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_1961_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_1961_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_1961_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_1961_inst_ack_1 : boolean;
  signal W_num_done_2169_delayed_2_0_2256_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_2191_inst_req_0 : boolean;
  signal W_read_k_2011_delayed_1_0_2073_inst_req_1 : boolean;
  signal type_cast_2262_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_1965_inst_req_0 : boolean;
  signal slice_2250_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_1965_inst_ack_0 : boolean;
  signal type_cast_2262_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_1965_inst_req_1 : boolean;
  signal slice_2250_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_1965_inst_ack_1 : boolean;
  signal W_num_done_2169_delayed_2_0_2256_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2260_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_1969_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_1969_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_1969_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_1969_inst_ack_1 : boolean;
  signal W_read_ip_1927_delayed_1_0_1971_inst_req_0 : boolean;
  signal W_read_ip_1927_delayed_1_0_1971_inst_ack_0 : boolean;
  signal W_read_ip_1927_delayed_1_0_1971_inst_req_1 : boolean;
  signal W_read_ip_1927_delayed_1_0_1971_inst_ack_1 : boolean;
  signal W_num_done_2169_delayed_2_0_2256_inst_ack_0 : boolean;
  signal W_store_kernel_2109_delayed_1_0_2187_inst_ack_1 : boolean;
  signal W_read_ip_1933_delayed_1_0_1980_inst_req_0 : boolean;
  signal W_read_ip_1933_delayed_1_0_1980_inst_ack_0 : boolean;
  signal W_read_ip_1933_delayed_1_0_1980_inst_req_1 : boolean;
  signal W_read_ip_1933_delayed_1_0_1980_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2260_inst_ack_1 : boolean;
  signal type_cast_2270_inst_req_1 : boolean;
  signal W_store_kernel_2109_delayed_1_0_2187_inst_req_1 : boolean;
  signal W_read_ip_1939_delayed_1_0_1989_inst_req_0 : boolean;
  signal W_num_done_2156_delayed_1_0_2239_inst_ack_1 : boolean;
  signal W_read_ip_1939_delayed_1_0_1989_inst_ack_0 : boolean;
  signal W_read_ip_1939_delayed_1_0_1989_inst_req_1 : boolean;
  signal W_num_done_2156_delayed_1_0_2239_inst_req_1 : boolean;
  signal W_read_ip_1939_delayed_1_0_1989_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_2260_inst_req_1 : boolean;
  signal type_cast_2270_inst_req_0 : boolean;
  signal W_num_done_2174_delayed_2_0_2264_inst_ack_0 : boolean;
  signal W_store_kernel_2109_delayed_1_0_2187_inst_ack_0 : boolean;
  signal W_write_input_1953_delayed_1_0_2007_inst_req_0 : boolean;
  signal W_write_input_1953_delayed_1_0_2007_inst_ack_0 : boolean;
  signal W_write_input_1953_delayed_1_0_2007_inst_req_1 : boolean;
  signal W_write_input_1953_delayed_1_0_2007_inst_ack_1 : boolean;
  signal W_num_done_2156_delayed_1_0_2239_inst_ack_0 : boolean;
  signal W_read_k_2023_delayed_1_0_2091_inst_ack_1 : boolean;
  signal W_store_kernel_2109_delayed_1_0_2187_inst_req_0 : boolean;
  signal W_read_k_2023_delayed_1_0_2091_inst_req_1 : boolean;
  signal type_cast_2262_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2011_inst_req_0 : boolean;
  signal W_num_done_2156_delayed_1_0_2239_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2011_inst_ack_0 : boolean;
  signal type_cast_2262_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2011_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2011_inst_ack_1 : boolean;
  signal W_num_done_2169_delayed_2_0_2256_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_2184_inst_ack_1 : boolean;
  signal W_read_k_2011_delayed_1_0_2073_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_2184_inst_req_1 : boolean;
  signal W_write_input_1957_delayed_1_0_2014_inst_req_0 : boolean;
  signal W_write_input_1957_delayed_1_0_2014_inst_ack_0 : boolean;
  signal W_write_input_1957_delayed_1_0_2014_inst_req_1 : boolean;
  signal W_write_input_1957_delayed_1_0_2014_inst_ack_1 : boolean;
  signal W_read_k_2023_delayed_1_0_2091_inst_ack_0 : boolean;
  signal W_read_k_2023_delayed_1_0_2091_inst_req_0 : boolean;
  signal W_read_k_2011_delayed_1_0_2073_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_2184_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2018_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_2198_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2018_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2018_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2018_inst_ack_1 : boolean;
  signal W_write_input_1961_delayed_1_0_2021_inst_req_0 : boolean;
  signal W_write_input_1961_delayed_1_0_2021_inst_ack_0 : boolean;
  signal W_write_input_1961_delayed_1_0_2021_inst_req_1 : boolean;
  signal W_write_input_1961_delayed_1_0_2021_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2025_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2025_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2025_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2025_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe1_2051_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe1_2051_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe1_2051_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe1_2051_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe2_2055_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe2_2055_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe2_2055_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe2_2055_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe3_2059_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe3_2059_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe3_2059_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe3_2059_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2063_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2063_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2063_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2063_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2067_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2067_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2067_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2067_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2071_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2071_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2071_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2071_inst_ack_1 : boolean;
  signal do_while_stmt_1908_branch_ack_0 : boolean;
  signal do_while_stmt_1908_branch_ack_1 : boolean;
  signal WPIPE_input_done_pipe_2275_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_2275_inst_ack_0 : boolean;
  signal WPIPE_input_done_pipe_2275_inst_req_1 : boolean;
  signal WPIPE_input_done_pipe_2275_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolve_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolve_CP_4643_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolve_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_4643_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolve_CP_4643_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_4643_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolve_CP_4643: Block -- control-path 
    signal convolve_CP_4643_elements: BooleanArray(281 downto 0);
    -- 
  begin -- 
    convolve_CP_4643_elements(0) <= convolve_CP_4643_start;
    convolve_CP_4643_symbol <= convolve_CP_4643_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	281 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1891/$entry
      -- CP-element group 0: 	 branch_block_stmt_1891/branch_block_stmt_1891__entry__
      -- CP-element group 0: 	 branch_block_stmt_1891/merge_stmt_1892__entry__
      -- CP-element group 0: 	 branch_block_stmt_1891/merge_stmt_1892_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1891/merge_stmt_1892__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_1891/merge_stmt_1892__entry___PhiReq/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1891/$exit
      -- CP-element group 1: 	 branch_block_stmt_1891/branch_block_stmt_1891__exit__
      -- 
    convolve_CP_4643_elements(1) <= false; 
    -- CP-element group 2:  transition  place  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	278 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	279 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1891/do_while_stmt_1908__exit__
      -- CP-element group 2: 	 branch_block_stmt_1891/assign_stmt_2277__entry__
      -- CP-element group 2: 	 branch_block_stmt_1891/assign_stmt_2277/$entry
      -- CP-element group 2: 	 branch_block_stmt_1891/assign_stmt_2277/WPIPE_input_done_pipe_2275_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1891/assign_stmt_2277/WPIPE_input_done_pipe_2275_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1891/assign_stmt_2277/WPIPE_input_done_pipe_2275_Sample/req
      -- 
    req_5567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(2), ack => WPIPE_input_done_pipe_2275_inst_req_0); -- 
    convolve_CP_4643_elements(2) <= convolve_CP_4643_elements(278);
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	281 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1894_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1894_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1894_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1894_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1894_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1894_Update/cr
      -- 
    ra_4675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1894_inst_ack_0, ack => convolve_CP_4643_elements(3)); -- 
    cr_4679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(3), ack => RPIPE_num_out_pipe_1894_inst_req_1); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1896_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1894_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1894_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1894_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1896_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1896_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1899_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1899_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1899_Sample/rr
      -- 
    ca_4680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1894_inst_ack_1, ack => convolve_CP_4643_elements(4)); -- 
    rr_4684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(4), ack => SUB_u16_u16_1896_inst_req_0); -- 
    rr_4702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(4), ack => RPIPE_num_out_pipe_1899_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1896_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1896_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1896_Sample/ra
      -- 
    ra_4685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_1896_inst_ack_0, ack => convolve_CP_4643_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	281 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	15 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1896_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1896_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1896_Update/ca
      -- 
    ca_4690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_1896_inst_ack_1, ack => convolve_CP_4643_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1899_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1899_update_start_
      -- CP-element group 7: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1899_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1899_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1899_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1899_Update/cr
      -- 
    ra_4703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1899_inst_ack_0, ack => convolve_CP_4643_elements(7)); -- 
    cr_4707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(7), ack => RPIPE_num_out_pipe_1899_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1901_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1899_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1899_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1899_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1901_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1901_Sample/rr
      -- 
    ca_4708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1899_inst_ack_1, ack => convolve_CP_4643_elements(8)); -- 
    rr_4712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(8), ack => SUB_u16_u16_1901_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1901_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1901_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1901_Sample/ra
      -- 
    ra_4713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_1901_inst_ack_0, ack => convolve_CP_4643_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	281 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	15 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1901_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1901_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1901_Update/ca
      -- 
    ca_4718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_1901_inst_ack_1, ack => convolve_CP_4643_elements(10)); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	281 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_size_pipe_1904_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_size_pipe_1904_update_start_
      -- CP-element group 11: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_size_pipe_1904_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_size_pipe_1904_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_size_pipe_1904_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_size_pipe_1904_Update/cr
      -- 
    ra_4731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1904_inst_ack_0, ack => convolve_CP_4643_elements(11)); -- 
    cr_4735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(11), ack => RPIPE_size_pipe_1904_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1906_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_size_pipe_1904_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_size_pipe_1904_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_size_pipe_1904_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1906_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1906_Sample/rr
      -- 
    ca_4736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1904_inst_ack_1, ack => convolve_CP_4643_elements(12)); -- 
    rr_4740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(12), ack => SUB_u16_u16_1906_inst_req_0); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1906_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1906_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1906_Sample/ra
      -- 
    ra_4741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_1906_inst_ack_0, ack => convolve_CP_4643_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	281 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1906_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1906_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1906_Update/ca
      -- 
    ca_4746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_1906_inst_ack_1, ack => convolve_CP_4643_elements(14)); -- 
    -- CP-element group 15:  join  transition  place  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	6 
    -- CP-element group 15: 	10 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907__exit__
      -- CP-element group 15: 	 branch_block_stmt_1891/do_while_stmt_1908__entry__
      -- CP-element group 15: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/$exit
      -- 
    convolve_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(6) & convolve_CP_4643_elements(10) & convolve_CP_4643_elements(14);
      gj_convolve_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  transition  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	22 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_1891/do_while_stmt_1908/$entry
      -- CP-element group 16: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908__entry__
      -- 
    convolve_CP_4643_elements(16) <= convolve_CP_4643_elements(15);
    -- CP-element group 17:  merge  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	278 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908__exit__
      -- 
    -- Element group convolve_CP_4643_elements(17) is bound as output of CP function.
    -- CP-element group 18:  merge  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1891/do_while_stmt_1908/loop_back
      -- 
    -- Element group convolve_CP_4643_elements(18) is bound as output of CP function.
    -- CP-element group 19:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	24 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	276 
    -- CP-element group 19: 	277 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1891/do_while_stmt_1908/condition_done
      -- CP-element group 19: 	 branch_block_stmt_1891/do_while_stmt_1908/loop_exit/$entry
      -- CP-element group 19: 	 branch_block_stmt_1891/do_while_stmt_1908/loop_taken/$entry
      -- 
    convolve_CP_4643_elements(19) <= convolve_CP_4643_elements(24);
    -- CP-element group 20:  branch  place  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	275 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1891/do_while_stmt_1908/loop_body_done
      -- 
    convolve_CP_4643_elements(20) <= convolve_CP_4643_elements(275);
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	33 
    -- CP-element group 21: 	90 
    -- CP-element group 21: 	109 
    -- CP-element group 21: 	71 
    -- CP-element group 21: 	52 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/back_edge_to_loop_body
      -- 
    convolve_CP_4643_elements(21) <= convolve_CP_4643_elements(18);
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	16 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	73 
    -- CP-element group 22: 	92 
    -- CP-element group 22: 	111 
    -- CP-element group 22: 	54 
    -- CP-element group 22: 	35 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/first_time_through_loop_body
      -- 
    convolve_CP_4643_elements(22) <= convolve_CP_4643_elements(16);
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	29 
    -- CP-element group 23: 	30 
    -- CP-element group 23: 	84 
    -- CP-element group 23: 	85 
    -- CP-element group 23: 	122 
    -- CP-element group 23: 	103 
    -- CP-element group 23: 	104 
    -- CP-element group 23: 	126 
    -- CP-element group 23: 	130 
    -- CP-element group 23: 	134 
    -- CP-element group 23: 	138 
    -- CP-element group 23: 	65 
    -- CP-element group 23: 	66 
    -- CP-element group 23: 	142 
    -- CP-element group 23: 	191 
    -- CP-element group 23: 	195 
    -- CP-element group 23: 	199 
    -- CP-element group 23: 	46 
    -- CP-element group 23: 	47 
    -- CP-element group 23: 	183 
    -- CP-element group 23: 	187 
    -- CP-element group 23: 	179 
    -- CP-element group 23: 	274 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/loop_body_start
      -- CP-element group 23: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/$entry
      -- 
    -- Element group convolve_CP_4643_elements(23) is bound as output of CP function.
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	89 
    -- CP-element group 24: 	108 
    -- CP-element group 24: 	70 
    -- CP-element group 24: 	51 
    -- CP-element group 24: 	274 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	19 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/condition_evaluated
      -- 
    condition_evaluated_4761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_4761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(24), ack => do_while_stmt_1908_branch_req_0); -- 
    convolve_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(28) & convolve_CP_4643_elements(89) & convolve_CP_4643_elements(108) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(51) & convolve_CP_4643_elements(274);
      gj_convolve_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	29 
    -- CP-element group 25: 	84 
    -- CP-element group 25: 	103 
    -- CP-element group 25: 	65 
    -- CP-element group 25: 	46 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	28 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	86 
    -- CP-element group 25: 	105 
    -- CP-element group 25: 	67 
    -- CP-element group 25: 	48 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/aggregated_phi_sample_req
      -- CP-element group 25: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1910_sample_start__ps
      -- 
    convolve_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(29) & convolve_CP_4643_elements(84) & convolve_CP_4643_elements(103) & convolve_CP_4643_elements(65) & convolve_CP_4643_elements(46) & convolve_CP_4643_elements(28);
      gj_convolve_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	31 
    -- CP-element group 26: 	87 
    -- CP-element group 26: 	106 
    -- CP-element group 26: 	68 
    -- CP-element group 26: 	49 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	123 
    -- CP-element group 26: 	127 
    -- CP-element group 26: 	131 
    -- CP-element group 26: 	135 
    -- CP-element group 26: 	139 
    -- CP-element group 26: 	143 
    -- CP-element group 26: 	192 
    -- CP-element group 26: 	196 
    -- CP-element group 26: 	200 
    -- CP-element group 26: 	147 
    -- CP-element group 26: 	151 
    -- CP-element group 26: 	155 
    -- CP-element group 26: 	184 
    -- CP-element group 26: 	188 
    -- CP-element group 26: 	204 
    -- CP-element group 26: 	208 
    -- CP-element group 26: 	212 
    -- CP-element group 26: 	180 
    -- CP-element group 26: 	241 
    -- CP-element group 26: 	216 
    -- CP-element group 26: 	275 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	29 
    -- CP-element group 26: 	84 
    -- CP-element group 26: 	103 
    -- CP-element group 26: 	65 
    -- CP-element group 26: 	46 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1921_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/aggregated_phi_sample_ack
      -- CP-element group 26: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1910_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1926_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1916_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1932_sample_completed_
      -- 
    convolve_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(31) & convolve_CP_4643_elements(87) & convolve_CP_4643_elements(106) & convolve_CP_4643_elements(68) & convolve_CP_4643_elements(49);
      gj_convolve_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	30 
    -- CP-element group 27: 	85 
    -- CP-element group 27: 	104 
    -- CP-element group 27: 	66 
    -- CP-element group 27: 	47 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	88 
    -- CP-element group 27: 	107 
    -- CP-element group 27: 	69 
    -- CP-element group 27: 	50 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1910_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/aggregated_phi_update_req
      -- 
    convolve_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(30) & convolve_CP_4643_elements(85) & convolve_CP_4643_elements(104) & convolve_CP_4643_elements(66) & convolve_CP_4643_elements(47);
      gj_convolve_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	32 
    -- CP-element group 28: 	89 
    -- CP-element group 28: 	108 
    -- CP-element group 28: 	70 
    -- CP-element group 28: 	51 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	25 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/aggregated_phi_update_ack
      -- 
    convolve_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(32) & convolve_CP_4643_elements(89) & convolve_CP_4643_elements(108) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(51);
      gj_convolve_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	23 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: 	125 
    -- CP-element group 29: 	129 
    -- CP-element group 29: 	133 
    -- CP-element group 29: 	137 
    -- CP-element group 29: 	141 
    -- CP-element group 29: 	190 
    -- CP-element group 29: 	194 
    -- CP-element group 29: 	198 
    -- CP-element group 29: 	145 
    -- CP-element group 29: 	149 
    -- CP-element group 29: 	153 
    -- CP-element group 29: 	157 
    -- CP-element group 29: 	182 
    -- CP-element group 29: 	186 
    -- CP-element group 29: 	202 
    -- CP-element group 29: 	206 
    -- CP-element group 29: 	210 
    -- CP-element group 29: 	214 
    -- CP-element group 29: 	243 
    -- CP-element group 29: 	218 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	25 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1910_sample_start_
      -- 
    convolve_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 21) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_markings: IntegerArray(0 to 21)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1);
      constant place_delays: IntegerArray(0 to 21) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 22); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(26) & convolve_CP_4643_elements(125) & convolve_CP_4643_elements(129) & convolve_CP_4643_elements(133) & convolve_CP_4643_elements(137) & convolve_CP_4643_elements(141) & convolve_CP_4643_elements(190) & convolve_CP_4643_elements(194) & convolve_CP_4643_elements(198) & convolve_CP_4643_elements(145) & convolve_CP_4643_elements(149) & convolve_CP_4643_elements(153) & convolve_CP_4643_elements(157) & convolve_CP_4643_elements(182) & convolve_CP_4643_elements(186) & convolve_CP_4643_elements(202) & convolve_CP_4643_elements(206) & convolve_CP_4643_elements(210) & convolve_CP_4643_elements(214) & convolve_CP_4643_elements(243) & convolve_CP_4643_elements(218);
      gj_convolve_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 22, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	23 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: 	217 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	27 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1910_update_start_
      -- 
    convolve_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(32) & convolve_CP_4643_elements(217);
      gj_convolve_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	26 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1910_sample_completed__ps
      -- 
    -- Element group convolve_CP_4643_elements(31) is bound as output of CP function.
    -- CP-element group 32:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	28 
    -- CP-element group 32: 	215 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1910_update_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1910_update_completed_
      -- 
    -- Element group convolve_CP_4643_elements(32) is bound as output of CP function.
    -- CP-element group 33:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	21 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1910_loopback_trigger
      -- 
    convolve_CP_4643_elements(33) <= convolve_CP_4643_elements(21);
    -- CP-element group 34:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1910_loopback_sample_req_ps
      -- CP-element group 34: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1910_loopback_sample_req
      -- 
    phi_stmt_1910_loopback_sample_req_4776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1910_loopback_sample_req_4776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(34), ack => phi_stmt_1910_req_1); -- 
    -- Element group convolve_CP_4643_elements(34) is bound as output of CP function.
    -- CP-element group 35:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	22 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1910_entry_trigger
      -- 
    convolve_CP_4643_elements(35) <= convolve_CP_4643_elements(22);
    -- CP-element group 36:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (2) 
      -- CP-element group 36: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1910_entry_sample_req
      -- CP-element group 36: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1910_entry_sample_req_ps
      -- 
    phi_stmt_1910_entry_sample_req_4779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1910_entry_sample_req_4779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(36), ack => phi_stmt_1910_req_0); -- 
    -- Element group convolve_CP_4643_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1910_phi_mux_ack
      -- CP-element group 37: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1910_phi_mux_ack_ps
      -- 
    phi_stmt_1910_phi_mux_ack_4782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1910_ack_0, ack => convolve_CP_4643_elements(37)); -- 
    -- CP-element group 38:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1914_sample_start__ps
      -- CP-element group 38: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1914_sample_completed__ps
      -- CP-element group 38: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1914_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1914_sample_completed_
      -- 
    -- Element group convolve_CP_4643_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1914_update_start__ps
      -- CP-element group 39: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1914_update_start_
      -- 
    -- Element group convolve_CP_4643_elements(39) is bound as output of CP function.
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	41 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1914_update_completed__ps
      -- 
    convolve_CP_4643_elements(40) <= convolve_CP_4643_elements(41);
    -- CP-element group 41:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	40 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1914_update_completed_
      -- 
    -- Element group convolve_CP_4643_elements(41) is a control-delay.
    cp_element_41_delay: control_delay_element  generic map(name => " 41_delay", delay_value => 1)  port map(req => convolve_CP_4643_elements(39), ack => convolve_CP_4643_elements(41), clk => clk, reset =>reset);
    -- CP-element group 42:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (4) 
      -- CP-element group 42: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_nacc_1915_sample_start__ps
      -- CP-element group 42: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_nacc_1915_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_nacc_1915_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_nacc_1915_Sample/req
      -- 
    req_4803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(42), ack => nacc_2247_1915_buf_req_0); -- 
    -- Element group convolve_CP_4643_elements(42) is bound as output of CP function.
    -- CP-element group 43:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_nacc_1915_update_start_
      -- CP-element group 43: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_nacc_1915_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_nacc_1915_Update/req
      -- CP-element group 43: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_nacc_1915_update_start__ps
      -- 
    req_4808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(43), ack => nacc_2247_1915_buf_req_1); -- 
    -- Element group convolve_CP_4643_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (4) 
      -- CP-element group 44: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_nacc_1915_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_nacc_1915_sample_completed__ps
      -- CP-element group 44: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_nacc_1915_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_nacc_1915_Sample/ack
      -- 
    ack_4804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_2247_1915_buf_ack_0, ack => convolve_CP_4643_elements(44)); -- 
    -- CP-element group 45:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_nacc_1915_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_nacc_1915_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_nacc_1915_Update/ack
      -- CP-element group 45: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_nacc_1915_update_completed__ps
      -- 
    ack_4809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_2247_1915_buf_ack_1, ack => convolve_CP_4643_elements(45)); -- 
    -- CP-element group 46:  join  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	23 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	26 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	25 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1916_sample_start_
      -- 
    convolve_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(26);
      gj_convolve_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	23 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	192 
    -- CP-element group 47: 	196 
    -- CP-element group 47: 	200 
    -- CP-element group 47: 	51 
    -- CP-element group 47: 	228 
    -- CP-element group 47: 	184 
    -- CP-element group 47: 	188 
    -- CP-element group 47: 	205 
    -- CP-element group 47: 	209 
    -- CP-element group 47: 	213 
    -- CP-element group 47: 	180 
    -- CP-element group 47: 	235 
    -- CP-element group 47: 	221 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	27 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1916_update_start_
      -- 
    convolve_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(192) & convolve_CP_4643_elements(196) & convolve_CP_4643_elements(200) & convolve_CP_4643_elements(51) & convolve_CP_4643_elements(228) & convolve_CP_4643_elements(184) & convolve_CP_4643_elements(188) & convolve_CP_4643_elements(205) & convolve_CP_4643_elements(209) & convolve_CP_4643_elements(213) & convolve_CP_4643_elements(180) & convolve_CP_4643_elements(235) & convolve_CP_4643_elements(221);
      gj_convolve_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	25 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1916_sample_start__ps
      -- 
    convolve_CP_4643_elements(48) <= convolve_CP_4643_elements(25);
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	26 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1916_sample_completed__ps
      -- 
    -- Element group convolve_CP_4643_elements(49) is bound as output of CP function.
    -- CP-element group 50:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	27 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1916_update_start__ps
      -- 
    convolve_CP_4643_elements(50) <= convolve_CP_4643_elements(27);
    -- CP-element group 51:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	24 
    -- CP-element group 51: 	28 
    -- CP-element group 51: 	192 
    -- CP-element group 51: 	196 
    -- CP-element group 51: 	200 
    -- CP-element group 51: 	226 
    -- CP-element group 51: 	233 
    -- CP-element group 51: 	184 
    -- CP-element group 51: 	188 
    -- CP-element group 51: 	203 
    -- CP-element group 51: 	207 
    -- CP-element group 51: 	211 
    -- CP-element group 51: 	180 
    -- CP-element group 51: 	219 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	47 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1916_update_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1916_update_completed_
      -- 
    -- Element group convolve_CP_4643_elements(51) is bound as output of CP function.
    -- CP-element group 52:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	21 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1916_loopback_trigger
      -- 
    convolve_CP_4643_elements(52) <= convolve_CP_4643_elements(21);
    -- CP-element group 53:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1916_loopback_sample_req
      -- CP-element group 53: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1916_loopback_sample_req_ps
      -- 
    phi_stmt_1916_loopback_sample_req_4820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1916_loopback_sample_req_4820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(53), ack => phi_stmt_1916_req_1); -- 
    -- Element group convolve_CP_4643_elements(53) is bound as output of CP function.
    -- CP-element group 54:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	22 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1916_entry_trigger
      -- 
    convolve_CP_4643_elements(54) <= convolve_CP_4643_elements(22);
    -- CP-element group 55:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1916_entry_sample_req
      -- CP-element group 55: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1916_entry_sample_req_ps
      -- 
    phi_stmt_1916_entry_sample_req_4823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1916_entry_sample_req_4823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(55), ack => phi_stmt_1916_req_0); -- 
    -- Element group convolve_CP_4643_elements(55) is bound as output of CP function.
    -- CP-element group 56:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1916_phi_mux_ack
      -- CP-element group 56: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1916_phi_mux_ack_ps
      -- 
    phi_stmt_1916_phi_mux_ack_4826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1916_ack_0, ack => convolve_CP_4643_elements(56)); -- 
    -- CP-element group 57:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1919_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1919_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1919_sample_start__ps
      -- CP-element group 57: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1919_sample_completed__ps
      -- 
    -- Element group convolve_CP_4643_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1919_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1919_update_start__ps
      -- 
    -- Element group convolve_CP_4643_elements(58) is bound as output of CP function.
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1919_update_completed__ps
      -- 
    convolve_CP_4643_elements(59) <= convolve_CP_4643_elements(60);
    -- CP-element group 60:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	59 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1919_update_completed_
      -- 
    -- Element group convolve_CP_4643_elements(60) is a control-delay.
    cp_element_60_delay: control_delay_element  generic map(name => " 60_delay", delay_value => 1)  port map(req => convolve_CP_4643_elements(58), ack => convolve_CP_4643_elements(60), clk => clk, reset =>reset);
    -- CP-element group 61:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (4) 
      -- CP-element group 61: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_row_1920_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_row_1920_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_row_1920_sample_start__ps
      -- CP-element group 61: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_row_1920_Sample/req
      -- 
    req_4847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(61), ack => n_row_2238_1920_buf_req_0); -- 
    -- Element group convolve_CP_4643_elements(61) is bound as output of CP function.
    -- CP-element group 62:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_row_1920_update_start_
      -- CP-element group 62: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_row_1920_Update/req
      -- CP-element group 62: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_row_1920_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_row_1920_update_start__ps
      -- 
    req_4852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(62), ack => n_row_2238_1920_buf_req_1); -- 
    -- Element group convolve_CP_4643_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (4) 
      -- CP-element group 63: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_row_1920_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_row_1920_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_row_1920_sample_completed__ps
      -- CP-element group 63: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_row_1920_Sample/ack
      -- 
    ack_4848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_2238_1920_buf_ack_0, ack => convolve_CP_4643_elements(63)); -- 
    -- CP-element group 64:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_row_1920_Update/ack
      -- CP-element group 64: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_row_1920_update_completed__ps
      -- CP-element group 64: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_row_1920_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_row_1920_update_completed_
      -- 
    ack_4853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_2238_1920_buf_ack_1, ack => convolve_CP_4643_elements(64)); -- 
    -- CP-element group 65:  join  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	23 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	26 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	25 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1921_sample_start_
      -- 
    convolve_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(26);
      gj_convolve_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  join  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	23 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	123 
    -- CP-element group 66: 	127 
    -- CP-element group 66: 	131 
    -- CP-element group 66: 	135 
    -- CP-element group 66: 	70 
    -- CP-element group 66: 	139 
    -- CP-element group 66: 	143 
    -- CP-element group 66: 	192 
    -- CP-element group 66: 	196 
    -- CP-element group 66: 	200 
    -- CP-element group 66: 	148 
    -- CP-element group 66: 	152 
    -- CP-element group 66: 	156 
    -- CP-element group 66: 	167 
    -- CP-element group 66: 	174 
    -- CP-element group 66: 	160 
    -- CP-element group 66: 	228 
    -- CP-element group 66: 	184 
    -- CP-element group 66: 	188 
    -- CP-element group 66: 	205 
    -- CP-element group 66: 	209 
    -- CP-element group 66: 	213 
    -- CP-element group 66: 	180 
    -- CP-element group 66: 	235 
    -- CP-element group 66: 	221 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	27 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1921_update_start_
      -- 
    convolve_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 25) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1);
      constant place_markings: IntegerArray(0 to 25)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1);
      constant place_delays: IntegerArray(0 to 25) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 26); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(123) & convolve_CP_4643_elements(127) & convolve_CP_4643_elements(131) & convolve_CP_4643_elements(135) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(139) & convolve_CP_4643_elements(143) & convolve_CP_4643_elements(192) & convolve_CP_4643_elements(196) & convolve_CP_4643_elements(200) & convolve_CP_4643_elements(148) & convolve_CP_4643_elements(152) & convolve_CP_4643_elements(156) & convolve_CP_4643_elements(167) & convolve_CP_4643_elements(174) & convolve_CP_4643_elements(160) & convolve_CP_4643_elements(228) & convolve_CP_4643_elements(184) & convolve_CP_4643_elements(188) & convolve_CP_4643_elements(205) & convolve_CP_4643_elements(209) & convolve_CP_4643_elements(213) & convolve_CP_4643_elements(180) & convolve_CP_4643_elements(235) & convolve_CP_4643_elements(221);
      gj_convolve_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 26, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	25 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1921_sample_start__ps
      -- 
    convolve_CP_4643_elements(67) <= convolve_CP_4643_elements(25);
    -- CP-element group 68:  join  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	26 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1921_sample_completed__ps
      -- 
    -- Element group convolve_CP_4643_elements(68) is bound as output of CP function.
    -- CP-element group 69:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	27 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1921_update_start__ps
      -- 
    convolve_CP_4643_elements(69) <= convolve_CP_4643_elements(27);
    -- CP-element group 70:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	24 
    -- CP-element group 70: 	28 
    -- CP-element group 70: 	123 
    -- CP-element group 70: 	127 
    -- CP-element group 70: 	131 
    -- CP-element group 70: 	135 
    -- CP-element group 70: 	139 
    -- CP-element group 70: 	143 
    -- CP-element group 70: 	192 
    -- CP-element group 70: 	196 
    -- CP-element group 70: 	200 
    -- CP-element group 70: 	226 
    -- CP-element group 70: 	146 
    -- CP-element group 70: 	150 
    -- CP-element group 70: 	154 
    -- CP-element group 70: 	158 
    -- CP-element group 70: 	165 
    -- CP-element group 70: 	172 
    -- CP-element group 70: 	233 
    -- CP-element group 70: 	184 
    -- CP-element group 70: 	188 
    -- CP-element group 70: 	203 
    -- CP-element group 70: 	207 
    -- CP-element group 70: 	211 
    -- CP-element group 70: 	180 
    -- CP-element group 70: 	219 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	66 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1921_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1921_update_completed__ps
      -- 
    -- Element group convolve_CP_4643_elements(70) is bound as output of CP function.
    -- CP-element group 71:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	21 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1921_loopback_trigger
      -- 
    convolve_CP_4643_elements(71) <= convolve_CP_4643_elements(21);
    -- CP-element group 72:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1921_loopback_sample_req
      -- CP-element group 72: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1921_loopback_sample_req_ps
      -- 
    phi_stmt_1921_loopback_sample_req_4864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1921_loopback_sample_req_4864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(72), ack => phi_stmt_1921_req_1); -- 
    -- Element group convolve_CP_4643_elements(72) is bound as output of CP function.
    -- CP-element group 73:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	22 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1921_entry_trigger
      -- 
    convolve_CP_4643_elements(73) <= convolve_CP_4643_elements(22);
    -- CP-element group 74:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1921_entry_sample_req
      -- CP-element group 74: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1921_entry_sample_req_ps
      -- 
    phi_stmt_1921_entry_sample_req_4867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1921_entry_sample_req_4867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(74), ack => phi_stmt_1921_req_0); -- 
    -- Element group convolve_CP_4643_elements(74) is bound as output of CP function.
    -- CP-element group 75:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1921_phi_mux_ack
      -- CP-element group 75: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1921_phi_mux_ack_ps
      -- 
    phi_stmt_1921_phi_mux_ack_4870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1921_ack_0, ack => convolve_CP_4643_elements(75)); -- 
    -- CP-element group 76:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1924_sample_completed__ps
      -- CP-element group 76: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1924_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1924_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1924_sample_start__ps
      -- 
    -- Element group convolve_CP_4643_elements(76) is bound as output of CP function.
    -- CP-element group 77:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1924_update_start__ps
      -- CP-element group 77: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1924_update_start_
      -- 
    -- Element group convolve_CP_4643_elements(77) is bound as output of CP function.
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1924_update_completed__ps
      -- 
    convolve_CP_4643_elements(78) <= convolve_CP_4643_elements(79);
    -- CP-element group 79:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	78 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1924_update_completed_
      -- 
    -- Element group convolve_CP_4643_elements(79) is a control-delay.
    cp_element_79_delay: control_delay_element  generic map(name => " 79_delay", delay_value => 1)  port map(req => convolve_CP_4643_elements(77), ack => convolve_CP_4643_elements(79), clk => clk, reset =>reset);
    -- CP-element group 80:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_col_1925_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_col_1925_Sample/req
      -- CP-element group 80: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_col_1925_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_col_1925_sample_start__ps
      -- 
    req_4891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(80), ack => n_col_2230_1925_buf_req_0); -- 
    -- Element group convolve_CP_4643_elements(80) is bound as output of CP function.
    -- CP-element group 81:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_col_1925_Update/req
      -- CP-element group 81: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_col_1925_update_start_
      -- CP-element group 81: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_col_1925_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_col_1925_update_start__ps
      -- 
    req_4896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(81), ack => n_col_2230_1925_buf_req_1); -- 
    -- Element group convolve_CP_4643_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_col_1925_Sample/ack
      -- CP-element group 82: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_col_1925_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_col_1925_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_col_1925_sample_completed__ps
      -- 
    ack_4892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_2230_1925_buf_ack_0, ack => convolve_CP_4643_elements(82)); -- 
    -- CP-element group 83:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_col_1925_update_completed__ps
      -- CP-element group 83: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_col_1925_Update/ack
      -- CP-element group 83: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_col_1925_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_col_1925_update_completed_
      -- 
    ack_4897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_2230_1925_buf_ack_1, ack => convolve_CP_4643_elements(83)); -- 
    -- CP-element group 84:  join  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	23 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	26 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	25 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1926_sample_start_
      -- 
    convolve_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(26);
      gj_convolve_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	23 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	89 
    -- CP-element group 85: 	123 
    -- CP-element group 85: 	127 
    -- CP-element group 85: 	131 
    -- CP-element group 85: 	135 
    -- CP-element group 85: 	139 
    -- CP-element group 85: 	143 
    -- CP-element group 85: 	148 
    -- CP-element group 85: 	152 
    -- CP-element group 85: 	156 
    -- CP-element group 85: 	167 
    -- CP-element group 85: 	174 
    -- CP-element group 85: 	160 
    -- CP-element group 85: 	242 
    -- CP-element group 85: 	254 
    -- CP-element group 85: 	265 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	27 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1926_update_start_
      -- 
    convolve_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(89) & convolve_CP_4643_elements(123) & convolve_CP_4643_elements(127) & convolve_CP_4643_elements(131) & convolve_CP_4643_elements(135) & convolve_CP_4643_elements(139) & convolve_CP_4643_elements(143) & convolve_CP_4643_elements(148) & convolve_CP_4643_elements(152) & convolve_CP_4643_elements(156) & convolve_CP_4643_elements(167) & convolve_CP_4643_elements(174) & convolve_CP_4643_elements(160) & convolve_CP_4643_elements(242) & convolve_CP_4643_elements(254) & convolve_CP_4643_elements(265);
      gj_convolve_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	25 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1926_sample_start__ps
      -- 
    convolve_CP_4643_elements(86) <= convolve_CP_4643_elements(25);
    -- CP-element group 87:  join  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	26 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1926_sample_completed__ps
      -- 
    -- Element group convolve_CP_4643_elements(87) is bound as output of CP function.
    -- CP-element group 88:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	27 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1926_update_start__ps
      -- 
    convolve_CP_4643_elements(88) <= convolve_CP_4643_elements(27);
    -- CP-element group 89:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	24 
    -- CP-element group 89: 	28 
    -- CP-element group 89: 	123 
    -- CP-element group 89: 	127 
    -- CP-element group 89: 	131 
    -- CP-element group 89: 	135 
    -- CP-element group 89: 	139 
    -- CP-element group 89: 	143 
    -- CP-element group 89: 	146 
    -- CP-element group 89: 	150 
    -- CP-element group 89: 	154 
    -- CP-element group 89: 	158 
    -- CP-element group 89: 	165 
    -- CP-element group 89: 	172 
    -- CP-element group 89: 	240 
    -- CP-element group 89: 	252 
    -- CP-element group 89: 	263 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	85 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1926_update_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1926_update_completed_
      -- 
    -- Element group convolve_CP_4643_elements(89) is bound as output of CP function.
    -- CP-element group 90:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	21 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1926_loopback_trigger
      -- 
    convolve_CP_4643_elements(90) <= convolve_CP_4643_elements(21);
    -- CP-element group 91:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1926_loopback_sample_req
      -- CP-element group 91: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1926_loopback_sample_req_ps
      -- 
    phi_stmt_1926_loopback_sample_req_4908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1926_loopback_sample_req_4908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(91), ack => phi_stmt_1926_req_1); -- 
    -- Element group convolve_CP_4643_elements(91) is bound as output of CP function.
    -- CP-element group 92:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	22 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1926_entry_trigger
      -- 
    convolve_CP_4643_elements(92) <= convolve_CP_4643_elements(22);
    -- CP-element group 93:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1926_entry_sample_req
      -- CP-element group 93: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1926_entry_sample_req_ps
      -- 
    phi_stmt_1926_entry_sample_req_4911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1926_entry_sample_req_4911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(93), ack => phi_stmt_1926_req_0); -- 
    -- Element group convolve_CP_4643_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1926_phi_mux_ack
      -- CP-element group 94: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1926_phi_mux_ack_ps
      -- 
    phi_stmt_1926_phi_mux_ack_4914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1926_ack_0, ack => convolve_CP_4643_elements(94)); -- 
    -- CP-element group 95:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1930_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1930_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1930_sample_start__ps
      -- CP-element group 95: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1930_sample_completed__ps
      -- 
    -- Element group convolve_CP_4643_elements(95) is bound as output of CP function.
    -- CP-element group 96:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1930_update_start_
      -- CP-element group 96: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1930_update_start__ps
      -- 
    -- Element group convolve_CP_4643_elements(96) is bound as output of CP function.
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1930_update_completed__ps
      -- 
    convolve_CP_4643_elements(97) <= convolve_CP_4643_elements(98);
    -- CP-element group 98:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	97 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1930_update_completed_
      -- 
    -- Element group convolve_CP_4643_elements(98) is a control-delay.
    cp_element_98_delay: control_delay_element  generic map(name => " 98_delay", delay_value => 1)  port map(req => convolve_CP_4643_elements(96), ack => convolve_CP_4643_elements(98), clk => clk, reset =>reset);
    -- CP-element group 99:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (4) 
      -- CP-element group 99: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_num_1931_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_num_1931_Sample/req
      -- CP-element group 99: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_num_1931_sample_start__ps
      -- CP-element group 99: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_num_1931_sample_start_
      -- 
    req_4935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(99), ack => n_num_2219_1931_buf_req_0); -- 
    -- Element group convolve_CP_4643_elements(99) is bound as output of CP function.
    -- CP-element group 100:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (4) 
      -- CP-element group 100: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_num_1931_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_num_1931_update_start_
      -- CP-element group 100: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_num_1931_Update/req
      -- CP-element group 100: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_num_1931_update_start__ps
      -- 
    req_4940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(100), ack => n_num_2219_1931_buf_req_1); -- 
    -- Element group convolve_CP_4643_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_num_1931_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_num_1931_Sample/ack
      -- CP-element group 101: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_num_1931_sample_completed__ps
      -- CP-element group 101: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_num_1931_sample_completed_
      -- 
    ack_4936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_num_2219_1931_buf_ack_0, ack => convolve_CP_4643_elements(101)); -- 
    -- CP-element group 102:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (4) 
      -- CP-element group 102: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_num_1931_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_num_1931_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_num_1931_Update/ack
      -- CP-element group 102: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_num_1931_update_completed__ps
      -- 
    ack_4941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_num_2219_1931_buf_ack_1, ack => convolve_CP_4643_elements(102)); -- 
    -- CP-element group 103:  join  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	23 
    -- CP-element group 103: marked-predecessors 
    -- CP-element group 103: 	26 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	25 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1932_sample_start_
      -- 
    convolve_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(26);
      gj_convolve_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  join  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	23 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	108 
    -- CP-element group 104: 	242 
    -- CP-element group 104: 	254 
    -- CP-element group 104: 	265 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	27 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1932_update_start_
      -- 
    convolve_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(108) & convolve_CP_4643_elements(242) & convolve_CP_4643_elements(254) & convolve_CP_4643_elements(265);
      gj_convolve_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	25 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1932_sample_start__ps
      -- 
    convolve_CP_4643_elements(105) <= convolve_CP_4643_elements(25);
    -- CP-element group 106:  join  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	26 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1932_sample_completed__ps
      -- 
    -- Element group convolve_CP_4643_elements(106) is bound as output of CP function.
    -- CP-element group 107:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	27 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1932_update_start__ps
      -- 
    convolve_CP_4643_elements(107) <= convolve_CP_4643_elements(27);
    -- CP-element group 108:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	24 
    -- CP-element group 108: 	28 
    -- CP-element group 108: 	240 
    -- CP-element group 108: 	252 
    -- CP-element group 108: 	263 
    -- CP-element group 108: marked-successors 
    -- CP-element group 108: 	104 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1932_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1932_update_completed__ps
      -- 
    -- Element group convolve_CP_4643_elements(108) is bound as output of CP function.
    -- CP-element group 109:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	21 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1932_loopback_trigger
      -- 
    convolve_CP_4643_elements(109) <= convolve_CP_4643_elements(21);
    -- CP-element group 110:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1932_loopback_sample_req
      -- CP-element group 110: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1932_loopback_sample_req_ps
      -- 
    phi_stmt_1932_loopback_sample_req_4952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1932_loopback_sample_req_4952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(110), ack => phi_stmt_1932_req_1); -- 
    -- Element group convolve_CP_4643_elements(110) is bound as output of CP function.
    -- CP-element group 111:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	22 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1932_entry_trigger
      -- 
    convolve_CP_4643_elements(111) <= convolve_CP_4643_elements(22);
    -- CP-element group 112:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1932_entry_sample_req_ps
      -- CP-element group 112: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1932_entry_sample_req
      -- 
    phi_stmt_1932_entry_sample_req_4955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1932_entry_sample_req_4955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(112), ack => phi_stmt_1932_req_0); -- 
    -- Element group convolve_CP_4643_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1932_phi_mux_ack_ps
      -- CP-element group 113: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/phi_stmt_1932_phi_mux_ack
      -- 
    phi_stmt_1932_phi_mux_ack_4958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1932_ack_0, ack => convolve_CP_4643_elements(113)); -- 
    -- CP-element group 114:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1935_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1935_sample_start__ps
      -- CP-element group 114: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1935_sample_completed__ps
      -- CP-element group 114: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1935_sample_start_
      -- 
    -- Element group convolve_CP_4643_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1935_update_start_
      -- CP-element group 115: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1935_update_start__ps
      -- 
    -- Element group convolve_CP_4643_elements(115) is bound as output of CP function.
    -- CP-element group 116:  join  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1935_update_completed__ps
      -- 
    convolve_CP_4643_elements(116) <= convolve_CP_4643_elements(117);
    -- CP-element group 117:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	116 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_1935_update_completed_
      -- 
    -- Element group convolve_CP_4643_elements(117) is a control-delay.
    cp_element_117_delay: control_delay_element  generic map(name => " 117_delay", delay_value => 1)  port map(req => convolve_CP_4643_elements(115), ack => convolve_CP_4643_elements(117), clk => clk, reset =>reset);
    -- CP-element group 118:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (4) 
      -- CP-element group 118: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_chl_1936_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_chl_1936_Sample/req
      -- CP-element group 118: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_chl_1936_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_chl_1936_sample_start__ps
      -- 
    req_4979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(118), ack => n_chl_2208_1936_buf_req_0); -- 
    -- Element group convolve_CP_4643_elements(118) is bound as output of CP function.
    -- CP-element group 119:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (4) 
      -- CP-element group 119: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_chl_1936_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_chl_1936_update_start_
      -- CP-element group 119: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_chl_1936_update_start__ps
      -- CP-element group 119: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_chl_1936_Update/req
      -- 
    req_4984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(119), ack => n_chl_2208_1936_buf_req_1); -- 
    -- Element group convolve_CP_4643_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (4) 
      -- CP-element group 120: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_chl_1936_Sample/ack
      -- CP-element group 120: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_chl_1936_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_chl_1936_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_chl_1936_sample_completed__ps
      -- 
    ack_4980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_2208_1936_buf_ack_0, ack => convolve_CP_4643_elements(120)); -- 
    -- CP-element group 121:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (4) 
      -- CP-element group 121: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_chl_1936_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_chl_1936_update_completed__ps
      -- CP-element group 121: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_chl_1936_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/R_n_chl_1936_Update/ack
      -- 
    ack_4985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_2208_1936_buf_ack_1, ack => convolve_CP_4643_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	23 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	125 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe1_1949_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe1_1949_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe1_1949_Sample/rr
      -- 
    rr_4994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(122), ack => RPIPE_input_pipe1_1949_inst_req_0); -- 
    convolve_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(125);
      gj_convolve_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	26 
    -- CP-element group 123: 	89 
    -- CP-element group 123: 	124 
    -- CP-element group 123: 	70 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	163 
    -- CP-element group 123: 	246 
    -- CP-element group 123: 	250 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	85 
    -- CP-element group 123: 	66 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe1_1949_update_start_
      -- CP-element group 123: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe1_1949_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe1_1949_Update/cr
      -- 
    cr_4999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(123), ack => RPIPE_input_pipe1_1949_inst_req_1); -- 
    convolve_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 1,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(89) & convolve_CP_4643_elements(124) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(163) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250);
      gj_convolve_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	123 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe1_1949_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe1_1949_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe1_1949_Sample/ra
      -- 
    ra_4995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1949_inst_ack_0, ack => convolve_CP_4643_elements(124)); -- 
    -- CP-element group 125:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	162 
    -- CP-element group 125: 	244 
    -- CP-element group 125: 	248 
    -- CP-element group 125: marked-successors 
    -- CP-element group 125: 	29 
    -- CP-element group 125: 	122 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe1_1949_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe1_1949_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe1_1949_Update/ca
      -- 
    ca_5000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1949_inst_ack_1, ack => convolve_CP_4643_elements(125)); -- 
    -- CP-element group 126:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	23 
    -- CP-element group 126: marked-predecessors 
    -- CP-element group 126: 	129 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe2_1953_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe2_1953_Sample/$entry
      -- CP-element group 126: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe2_1953_Sample/rr
      -- 
    rr_5008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(126), ack => RPIPE_input_pipe2_1953_inst_req_0); -- 
    convolve_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(129);
      gj_convolve_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	26 
    -- CP-element group 127: 	89 
    -- CP-element group 127: 	128 
    -- CP-element group 127: 	70 
    -- CP-element group 127: marked-predecessors 
    -- CP-element group 127: 	170 
    -- CP-element group 127: 	246 
    -- CP-element group 127: 	250 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	85 
    -- CP-element group 127: 	66 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe2_1953_update_start_
      -- CP-element group 127: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe2_1953_Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe2_1953_Update/cr
      -- 
    cr_5013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(127), ack => RPIPE_input_pipe2_1953_inst_req_1); -- 
    convolve_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 1,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(89) & convolve_CP_4643_elements(128) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(170) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250);
      gj_convolve_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	127 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe2_1953_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe2_1953_Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe2_1953_Sample/ra
      -- 
    ra_5009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe2_1953_inst_ack_0, ack => convolve_CP_4643_elements(128)); -- 
    -- CP-element group 129:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	169 
    -- CP-element group 129: 	244 
    -- CP-element group 129: 	248 
    -- CP-element group 129: marked-successors 
    -- CP-element group 129: 	29 
    -- CP-element group 129: 	126 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe2_1953_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe2_1953_Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe2_1953_Update/ca
      -- 
    ca_5014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe2_1953_inst_ack_1, ack => convolve_CP_4643_elements(129)); -- 
    -- CP-element group 130:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	23 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	133 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe3_1957_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe3_1957_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe3_1957_Sample/rr
      -- 
    rr_5022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(130), ack => RPIPE_input_pipe3_1957_inst_req_0); -- 
    convolve_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(133);
      gj_convolve_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	26 
    -- CP-element group 131: 	89 
    -- CP-element group 131: 	132 
    -- CP-element group 131: 	70 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	177 
    -- CP-element group 131: 	246 
    -- CP-element group 131: 	250 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	85 
    -- CP-element group 131: 	66 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe3_1957_update_start_
      -- CP-element group 131: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe3_1957_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe3_1957_Update/cr
      -- 
    cr_5027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(131), ack => RPIPE_input_pipe3_1957_inst_req_1); -- 
    convolve_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 1,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(89) & convolve_CP_4643_elements(132) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(177) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250);
      gj_convolve_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	131 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe3_1957_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe3_1957_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe3_1957_Sample/ra
      -- 
    ra_5023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe3_1957_inst_ack_0, ack => convolve_CP_4643_elements(132)); -- 
    -- CP-element group 133:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	176 
    -- CP-element group 133: 	244 
    -- CP-element group 133: 	248 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	29 
    -- CP-element group 133: 	130 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe3_1957_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe3_1957_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_input_pipe3_1957_Update/ca
      -- 
    ca_5028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe3_1957_inst_ack_1, ack => convolve_CP_4643_elements(133)); -- 
    -- CP-element group 134:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	23 
    -- CP-element group 134: marked-predecessors 
    -- CP-element group 134: 	137 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip1_1961_sample_start_
      -- CP-element group 134: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip1_1961_Sample/$entry
      -- CP-element group 134: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip1_1961_Sample/rr
      -- 
    rr_5036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(134), ack => RPIPE_xxconvolvexxconv_ip1_1961_inst_req_0); -- 
    convolve_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(137);
      gj_convolve_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	26 
    -- CP-element group 135: 	89 
    -- CP-element group 135: 	136 
    -- CP-element group 135: 	70 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	163 
    -- CP-element group 135: 	246 
    -- CP-element group 135: 	250 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135: marked-successors 
    -- CP-element group 135: 	85 
    -- CP-element group 135: 	66 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip1_1961_update_start_
      -- CP-element group 135: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip1_1961_Update/$entry
      -- CP-element group 135: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip1_1961_Update/cr
      -- 
    cr_5041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(135), ack => RPIPE_xxconvolvexxconv_ip1_1961_inst_req_1); -- 
    convolve_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 1,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(89) & convolve_CP_4643_elements(136) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(163) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250);
      gj_convolve_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  transition  input  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	135 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip1_1961_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip1_1961_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip1_1961_Sample/ra
      -- 
    ra_5037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip1_1961_inst_ack_0, ack => convolve_CP_4643_elements(136)); -- 
    -- CP-element group 137:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	162 
    -- CP-element group 137: 	244 
    -- CP-element group 137: 	248 
    -- CP-element group 137: marked-successors 
    -- CP-element group 137: 	29 
    -- CP-element group 137: 	134 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip1_1961_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip1_1961_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip1_1961_Update/ca
      -- 
    ca_5042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip1_1961_inst_ack_1, ack => convolve_CP_4643_elements(137)); -- 
    -- CP-element group 138:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	23 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	141 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip2_1965_sample_start_
      -- CP-element group 138: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip2_1965_Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip2_1965_Sample/rr
      -- 
    rr_5050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(138), ack => RPIPE_xxconvolvexxconv_ip2_1965_inst_req_0); -- 
    convolve_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(141);
      gj_convolve_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	26 
    -- CP-element group 139: 	89 
    -- CP-element group 139: 	70 
    -- CP-element group 139: 	140 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	170 
    -- CP-element group 139: 	246 
    -- CP-element group 139: 	250 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	85 
    -- CP-element group 139: 	66 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip2_1965_update_start_
      -- CP-element group 139: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip2_1965_Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip2_1965_Update/cr
      -- 
    cr_5055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(139), ack => RPIPE_xxconvolvexxconv_ip2_1965_inst_req_1); -- 
    convolve_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(89) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(140) & convolve_CP_4643_elements(170) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250);
      gj_convolve_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	139 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip2_1965_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip2_1965_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip2_1965_Sample/ra
      -- 
    ra_5051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip2_1965_inst_ack_0, ack => convolve_CP_4643_elements(140)); -- 
    -- CP-element group 141:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	169 
    -- CP-element group 141: 	244 
    -- CP-element group 141: 	248 
    -- CP-element group 141: marked-successors 
    -- CP-element group 141: 	29 
    -- CP-element group 141: 	138 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip2_1965_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip2_1965_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip2_1965_Update/ca
      -- 
    ca_5056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip2_1965_inst_ack_1, ack => convolve_CP_4643_elements(141)); -- 
    -- CP-element group 142:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	23 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	145 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip3_1969_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip3_1969_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip3_1969_Sample/rr
      -- 
    rr_5064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(142), ack => RPIPE_xxconvolvexxconv_ip3_1969_inst_req_0); -- 
    convolve_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(145);
      gj_convolve_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	26 
    -- CP-element group 143: 	89 
    -- CP-element group 143: 	70 
    -- CP-element group 143: 	144 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	177 
    -- CP-element group 143: 	246 
    -- CP-element group 143: 	250 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143: marked-successors 
    -- CP-element group 143: 	85 
    -- CP-element group 143: 	66 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip3_1969_update_start_
      -- CP-element group 143: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip3_1969_Update/$entry
      -- CP-element group 143: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip3_1969_Update/cr
      -- 
    cr_5069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(143), ack => RPIPE_xxconvolvexxconv_ip3_1969_inst_req_1); -- 
    convolve_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(89) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(144) & convolve_CP_4643_elements(177) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250);
      gj_convolve_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	143 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip3_1969_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip3_1969_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip3_1969_Sample/ra
      -- 
    ra_5065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip3_1969_inst_ack_0, ack => convolve_CP_4643_elements(144)); -- 
    -- CP-element group 145:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	176 
    -- CP-element group 145: 	244 
    -- CP-element group 145: 	248 
    -- CP-element group 145: marked-successors 
    -- CP-element group 145: 	29 
    -- CP-element group 145: 	142 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip3_1969_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip3_1969_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_ip3_1969_Update/ca
      -- 
    ca_5070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip3_1969_inst_ack_1, ack => convolve_CP_4643_elements(145)); -- 
    -- CP-element group 146:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	89 
    -- CP-element group 146: 	70 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	148 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1973_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1973_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1973_Sample/req
      -- 
    req_5078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(146), ack => W_read_ip_1927_delayed_1_0_1971_inst_req_0); -- 
    convolve_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(89) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(148);
      gj_convolve_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	26 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	149 
    -- CP-element group 147: 	163 
    -- CP-element group 147: 	246 
    -- CP-element group 147: 	250 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1973_update_start_
      -- CP-element group 147: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1973_Update/$entry
      -- CP-element group 147: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1973_Update/req
      -- 
    req_5083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(147), ack => W_read_ip_1927_delayed_1_0_1971_inst_req_1); -- 
    convolve_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(149) & convolve_CP_4643_elements(163) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250);
      gj_convolve_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	85 
    -- CP-element group 148: 	66 
    -- CP-element group 148: 	146 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1973_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1973_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1973_Sample/ack
      -- 
    ack_5079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_1927_delayed_1_0_1971_inst_ack_0, ack => convolve_CP_4643_elements(148)); -- 
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	162 
    -- CP-element group 149: 	244 
    -- CP-element group 149: 	248 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	29 
    -- CP-element group 149: 	147 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1973_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1973_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1973_Update/ack
      -- 
    ack_5084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_1927_delayed_1_0_1971_inst_ack_1, ack => convolve_CP_4643_elements(149)); -- 
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	89 
    -- CP-element group 150: 	70 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1982_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1982_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1982_Sample/req
      -- 
    req_5092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(150), ack => W_read_ip_1933_delayed_1_0_1980_inst_req_0); -- 
    convolve_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(89) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(152);
      gj_convolve_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	26 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: 	170 
    -- CP-element group 151: 	246 
    -- CP-element group 151: 	250 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1982_update_start_
      -- CP-element group 151: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1982_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1982_Update/req
      -- 
    req_5097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(151), ack => W_read_ip_1933_delayed_1_0_1980_inst_req_1); -- 
    convolve_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(153) & convolve_CP_4643_elements(170) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250);
      gj_convolve_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	85 
    -- CP-element group 152: 	66 
    -- CP-element group 152: 	150 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1982_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1982_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1982_Sample/ack
      -- 
    ack_5093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_1933_delayed_1_0_1980_inst_ack_0, ack => convolve_CP_4643_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	169 
    -- CP-element group 153: 	244 
    -- CP-element group 153: 	248 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	29 
    -- CP-element group 153: 	151 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1982_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1982_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1982_Update/ack
      -- 
    ack_5098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_1933_delayed_1_0_1980_inst_ack_1, ack => convolve_CP_4643_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	89 
    -- CP-element group 154: 	70 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1991_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1991_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1991_Sample/req
      -- 
    req_5106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(154), ack => W_read_ip_1939_delayed_1_0_1989_inst_req_0); -- 
    convolve_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(89) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(156);
      gj_convolve_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	26 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: 	177 
    -- CP-element group 155: 	246 
    -- CP-element group 155: 	250 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1991_update_start_
      -- CP-element group 155: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1991_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1991_Update/req
      -- 
    req_5111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(155), ack => W_read_ip_1939_delayed_1_0_1989_inst_req_1); -- 
    convolve_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(157) & convolve_CP_4643_elements(177) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250);
      gj_convolve_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	85 
    -- CP-element group 156: 	66 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1991_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1991_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1991_Sample/ack
      -- 
    ack_5107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_1939_delayed_1_0_1989_inst_ack_0, ack => convolve_CP_4643_elements(156)); -- 
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	176 
    -- CP-element group 157: 	244 
    -- CP-element group 157: 	248 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	29 
    -- CP-element group 157: 	155 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1991_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1991_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_1991_Update/ack
      -- 
    ack_5112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_1939_delayed_1_0_1989_inst_ack_1, ack => convolve_CP_4643_elements(157)); -- 
    -- CP-element group 158:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	89 
    -- CP-element group 158: 	70 
    -- CP-element group 158: marked-predecessors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2009_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2009_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2009_Sample/req
      -- 
    req_5120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(158), ack => W_write_input_1953_delayed_1_0_2007_inst_req_0); -- 
    convolve_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(89) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(160);
      gj_convolve_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: 	163 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2009_update_start_
      -- CP-element group 159: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2009_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2009_Update/req
      -- 
    req_5125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(159), ack => W_write_input_1953_delayed_1_0_2007_inst_req_1); -- 
    convolve_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(161) & convolve_CP_4643_elements(163);
      gj_convolve_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	85 
    -- CP-element group 160: 	66 
    -- CP-element group 160: 	158 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2009_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2009_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2009_Sample/ack
      -- 
    ack_5121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_1953_delayed_1_0_2007_inst_ack_0, ack => convolve_CP_4643_elements(160)); -- 
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	159 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2009_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2009_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2009_Update/ack
      -- 
    ack_5126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_1953_delayed_1_0_2007_inst_ack_1, ack => convolve_CP_4643_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	125 
    -- CP-element group 162: 	137 
    -- CP-element group 162: 	149 
    -- CP-element group 162: 	161 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip1_2011_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip1_2011_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip1_2011_Sample/req
      -- 
    req_5134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(162), ack => WPIPE_xxconvolvexxconv_ip1_2011_inst_req_0); -- 
    convolve_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(125) & convolve_CP_4643_elements(137) & convolve_CP_4643_elements(149) & convolve_CP_4643_elements(161) & convolve_CP_4643_elements(164);
      gj_convolve_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163: marked-successors 
    -- CP-element group 163: 	123 
    -- CP-element group 163: 	135 
    -- CP-element group 163: 	147 
    -- CP-element group 163: 	159 
    -- CP-element group 163:  members (6) 
      -- CP-element group 163: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip1_2011_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip1_2011_update_start_
      -- CP-element group 163: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip1_2011_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip1_2011_Sample/ack
      -- CP-element group 163: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip1_2011_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip1_2011_Update/req
      -- 
    ack_5135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip1_2011_inst_ack_0, ack => convolve_CP_4643_elements(163)); -- 
    req_5139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(163), ack => WPIPE_xxconvolvexxconv_ip1_2011_inst_req_1); -- 
    -- CP-element group 164:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	275 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	162 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip1_2011_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip1_2011_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip1_2011_Update/ack
      -- 
    ack_5140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip1_2011_inst_ack_1, ack => convolve_CP_4643_elements(164)); -- 
    -- CP-element group 165:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	89 
    -- CP-element group 165: 	70 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	167 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2016_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2016_Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2016_Sample/req
      -- 
    req_5148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(165), ack => W_write_input_1957_delayed_1_0_2014_inst_req_0); -- 
    convolve_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(89) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(167);
      gj_convolve_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	168 
    -- CP-element group 166: 	170 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2016_update_start_
      -- CP-element group 166: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2016_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2016_Update/req
      -- 
    req_5153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(166), ack => W_write_input_1957_delayed_1_0_2014_inst_req_1); -- 
    convolve_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(168) & convolve_CP_4643_elements(170);
      gj_convolve_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: marked-successors 
    -- CP-element group 167: 	85 
    -- CP-element group 167: 	66 
    -- CP-element group 167: 	165 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2016_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2016_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2016_Sample/ack
      -- 
    ack_5149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_1957_delayed_1_0_2014_inst_ack_0, ack => convolve_CP_4643_elements(167)); -- 
    -- CP-element group 168:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168: marked-successors 
    -- CP-element group 168: 	166 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2016_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2016_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2016_Update/ack
      -- 
    ack_5154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_1957_delayed_1_0_2014_inst_ack_1, ack => convolve_CP_4643_elements(168)); -- 
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	129 
    -- CP-element group 169: 	141 
    -- CP-element group 169: 	153 
    -- CP-element group 169: 	168 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	171 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip2_2018_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip2_2018_Sample/$entry
      -- CP-element group 169: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip2_2018_Sample/req
      -- 
    req_5162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(169), ack => WPIPE_xxconvolvexxconv_ip2_2018_inst_req_0); -- 
    convolve_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(129) & convolve_CP_4643_elements(141) & convolve_CP_4643_elements(153) & convolve_CP_4643_elements(168) & convolve_CP_4643_elements(171);
      gj_convolve_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	127 
    -- CP-element group 170: 	139 
    -- CP-element group 170: 	151 
    -- CP-element group 170: 	166 
    -- CP-element group 170:  members (6) 
      -- CP-element group 170: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip2_2018_update_start_
      -- CP-element group 170: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip2_2018_sample_completed_
      -- CP-element group 170: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip2_2018_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip2_2018_Sample/ack
      -- CP-element group 170: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip2_2018_Update/$entry
      -- CP-element group 170: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip2_2018_Update/req
      -- 
    ack_5163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip2_2018_inst_ack_0, ack => convolve_CP_4643_elements(170)); -- 
    req_5167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(170), ack => WPIPE_xxconvolvexxconv_ip2_2018_inst_req_1); -- 
    -- CP-element group 171:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	275 
    -- CP-element group 171: marked-successors 
    -- CP-element group 171: 	169 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip2_2018_update_completed_
      -- CP-element group 171: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip2_2018_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip2_2018_Update/ack
      -- 
    ack_5168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip2_2018_inst_ack_1, ack => convolve_CP_4643_elements(171)); -- 
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	89 
    -- CP-element group 172: 	70 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	174 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2023_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2023_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2023_Sample/req
      -- 
    req_5176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(172), ack => W_write_input_1961_delayed_1_0_2021_inst_req_0); -- 
    convolve_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(89) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(174);
      gj_convolve_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: 	177 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2023_update_start_
      -- CP-element group 173: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2023_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2023_Update/req
      -- 
    req_5181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(173), ack => W_write_input_1961_delayed_1_0_2021_inst_req_1); -- 
    convolve_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(175) & convolve_CP_4643_elements(177);
      gj_convolve_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: marked-successors 
    -- CP-element group 174: 	85 
    -- CP-element group 174: 	66 
    -- CP-element group 174: 	172 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2023_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2023_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2023_Sample/ack
      -- 
    ack_5177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_1961_delayed_1_0_2021_inst_ack_0, ack => convolve_CP_4643_elements(174)); -- 
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2023_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2023_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2023_Update/ack
      -- 
    ack_5182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_1961_delayed_1_0_2021_inst_ack_1, ack => convolve_CP_4643_elements(175)); -- 
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	133 
    -- CP-element group 176: 	145 
    -- CP-element group 176: 	157 
    -- CP-element group 176: 	175 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	178 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip3_2025_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip3_2025_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip3_2025_Sample/req
      -- 
    req_5190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(176), ack => WPIPE_xxconvolvexxconv_ip3_2025_inst_req_0); -- 
    convolve_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(133) & convolve_CP_4643_elements(145) & convolve_CP_4643_elements(157) & convolve_CP_4643_elements(175) & convolve_CP_4643_elements(178);
      gj_convolve_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	131 
    -- CP-element group 177: 	143 
    -- CP-element group 177: 	155 
    -- CP-element group 177: 	173 
    -- CP-element group 177:  members (6) 
      -- CP-element group 177: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip3_2025_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip3_2025_update_start_
      -- CP-element group 177: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip3_2025_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip3_2025_Sample/ack
      -- CP-element group 177: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip3_2025_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip3_2025_Update/req
      -- 
    ack_5191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip3_2025_inst_ack_0, ack => convolve_CP_4643_elements(177)); -- 
    req_5195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(177), ack => WPIPE_xxconvolvexxconv_ip3_2025_inst_req_1); -- 
    -- CP-element group 178:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	275 
    -- CP-element group 178: marked-successors 
    -- CP-element group 178: 	176 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip3_2025_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip3_2025_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_ip3_2025_Update/ack
      -- 
    ack_5196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip3_2025_inst_ack_1, ack => convolve_CP_4643_elements(178)); -- 
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	23 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	182 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe1_2051_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe1_2051_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe1_2051_Sample/rr
      -- 
    rr_5204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(179), ack => RPIPE_kernel_pipe1_2051_inst_req_0); -- 
    convolve_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(182);
      gj_convolve_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	26 
    -- CP-element group 180: 	70 
    -- CP-element group 180: 	51 
    -- CP-element group 180: 	181 
    -- CP-element group 180: marked-predecessors 
    -- CP-element group 180: 	224 
    -- CP-element group 180: 	246 
    -- CP-element group 180: 	250 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	66 
    -- CP-element group 180: 	47 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe1_2051_update_start_
      -- CP-element group 180: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe1_2051_Update/$entry
      -- CP-element group 180: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe1_2051_Update/cr
      -- 
    cr_5209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(180), ack => RPIPE_kernel_pipe1_2051_inst_req_1); -- 
    convolve_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(51) & convolve_CP_4643_elements(181) & convolve_CP_4643_elements(224) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250);
      gj_convolve_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	180 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe1_2051_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe1_2051_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe1_2051_Sample/ra
      -- 
    ra_5205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_2051_inst_ack_0, ack => convolve_CP_4643_elements(181)); -- 
    -- CP-element group 182:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	223 
    -- CP-element group 182: 	244 
    -- CP-element group 182: 	248 
    -- CP-element group 182: marked-successors 
    -- CP-element group 182: 	29 
    -- CP-element group 182: 	179 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe1_2051_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe1_2051_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe1_2051_Update/ca
      -- 
    ca_5210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_2051_inst_ack_1, ack => convolve_CP_4643_elements(182)); -- 
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	23 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	186 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe2_2055_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe2_2055_Sample/$entry
      -- CP-element group 183: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe2_2055_Sample/rr
      -- 
    rr_5218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(183), ack => RPIPE_kernel_pipe2_2055_inst_req_0); -- 
    convolve_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(186);
      gj_convolve_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	26 
    -- CP-element group 184: 	70 
    -- CP-element group 184: 	51 
    -- CP-element group 184: 	185 
    -- CP-element group 184: marked-predecessors 
    -- CP-element group 184: 	231 
    -- CP-element group 184: 	246 
    -- CP-element group 184: 	250 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	66 
    -- CP-element group 184: 	47 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe2_2055_update_start_
      -- CP-element group 184: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe2_2055_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe2_2055_Update/cr
      -- 
    cr_5223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(184), ack => RPIPE_kernel_pipe2_2055_inst_req_1); -- 
    convolve_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(51) & convolve_CP_4643_elements(185) & convolve_CP_4643_elements(231) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250);
      gj_convolve_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	184 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe2_2055_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe2_2055_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe2_2055_Sample/ra
      -- 
    ra_5219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe2_2055_inst_ack_0, ack => convolve_CP_4643_elements(185)); -- 
    -- CP-element group 186:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	230 
    -- CP-element group 186: 	244 
    -- CP-element group 186: 	248 
    -- CP-element group 186: marked-successors 
    -- CP-element group 186: 	29 
    -- CP-element group 186: 	183 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe2_2055_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe2_2055_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe2_2055_Update/ca
      -- 
    ca_5224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe2_2055_inst_ack_1, ack => convolve_CP_4643_elements(186)); -- 
    -- CP-element group 187:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	23 
    -- CP-element group 187: marked-predecessors 
    -- CP-element group 187: 	190 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	189 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe3_2059_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe3_2059_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe3_2059_Sample/rr
      -- 
    rr_5232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(187), ack => RPIPE_kernel_pipe3_2059_inst_req_0); -- 
    convolve_cp_element_group_187: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_187"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(190);
      gj_convolve_cp_element_group_187 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(187), clk => clk, reset => reset); --
    end block;
    -- CP-element group 188:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	26 
    -- CP-element group 188: 	70 
    -- CP-element group 188: 	189 
    -- CP-element group 188: 	51 
    -- CP-element group 188: marked-predecessors 
    -- CP-element group 188: 	246 
    -- CP-element group 188: 	250 
    -- CP-element group 188: 	238 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	190 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	66 
    -- CP-element group 188: 	47 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe3_2059_update_start_
      -- CP-element group 188: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe3_2059_Update/$entry
      -- CP-element group 188: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe3_2059_Update/cr
      -- 
    cr_5237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(188), ack => RPIPE_kernel_pipe3_2059_inst_req_1); -- 
    convolve_cp_element_group_188: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 1,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_188"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(189) & convolve_CP_4643_elements(51) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250) & convolve_CP_4643_elements(238);
      gj_convolve_cp_element_group_188 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 189:  transition  input  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	187 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	188 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe3_2059_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe3_2059_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe3_2059_Sample/ra
      -- 
    ra_5233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe3_2059_inst_ack_0, ack => convolve_CP_4643_elements(189)); -- 
    -- CP-element group 190:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	244 
    -- CP-element group 190: 	248 
    -- CP-element group 190: 	237 
    -- CP-element group 190: marked-successors 
    -- CP-element group 190: 	29 
    -- CP-element group 190: 	187 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe3_2059_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe3_2059_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_kernel_pipe3_2059_Update/ca
      -- 
    ca_5238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe3_2059_inst_ack_1, ack => convolve_CP_4643_elements(190)); -- 
    -- CP-element group 191:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	23 
    -- CP-element group 191: marked-predecessors 
    -- CP-element group 191: 	194 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	193 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k1_2063_sample_start_
      -- CP-element group 191: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k1_2063_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k1_2063_Sample/rr
      -- 
    rr_5246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(191), ack => RPIPE_xxconvolvexxconv_k1_2063_inst_req_0); -- 
    convolve_cp_element_group_191: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_191"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(194);
      gj_convolve_cp_element_group_191 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 192:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	26 
    -- CP-element group 192: 	70 
    -- CP-element group 192: 	193 
    -- CP-element group 192: 	51 
    -- CP-element group 192: marked-predecessors 
    -- CP-element group 192: 	224 
    -- CP-element group 192: 	246 
    -- CP-element group 192: 	250 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	194 
    -- CP-element group 192: marked-successors 
    -- CP-element group 192: 	66 
    -- CP-element group 192: 	47 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k1_2063_update_start_
      -- CP-element group 192: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k1_2063_Update/$entry
      -- CP-element group 192: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k1_2063_Update/cr
      -- 
    cr_5251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(192), ack => RPIPE_xxconvolvexxconv_k1_2063_inst_req_1); -- 
    convolve_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 1,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(193) & convolve_CP_4643_elements(51) & convolve_CP_4643_elements(224) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250);
      gj_convolve_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  transition  input  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	191 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	192 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k1_2063_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k1_2063_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k1_2063_Sample/ra
      -- 
    ra_5247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k1_2063_inst_ack_0, ack => convolve_CP_4643_elements(193)); -- 
    -- CP-element group 194:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	192 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	223 
    -- CP-element group 194: 	244 
    -- CP-element group 194: 	248 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	29 
    -- CP-element group 194: 	191 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k1_2063_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k1_2063_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k1_2063_Update/ca
      -- 
    ca_5252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k1_2063_inst_ack_1, ack => convolve_CP_4643_elements(194)); -- 
    -- CP-element group 195:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	23 
    -- CP-element group 195: marked-predecessors 
    -- CP-element group 195: 	198 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	197 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k2_2067_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k2_2067_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k2_2067_Sample/rr
      -- 
    rr_5260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(195), ack => RPIPE_xxconvolvexxconv_k2_2067_inst_req_0); -- 
    convolve_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(198);
      gj_convolve_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	26 
    -- CP-element group 196: 	70 
    -- CP-element group 196: 	197 
    -- CP-element group 196: 	51 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	231 
    -- CP-element group 196: 	246 
    -- CP-element group 196: 	250 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: marked-successors 
    -- CP-element group 196: 	66 
    -- CP-element group 196: 	47 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k2_2067_update_start_
      -- CP-element group 196: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k2_2067_Update/$entry
      -- CP-element group 196: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k2_2067_Update/cr
      -- 
    cr_5265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(196), ack => RPIPE_xxconvolvexxconv_k2_2067_inst_req_1); -- 
    convolve_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 1,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(197) & convolve_CP_4643_elements(51) & convolve_CP_4643_elements(231) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250);
      gj_convolve_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  transition  input  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	195 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	196 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k2_2067_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k2_2067_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k2_2067_Sample/ra
      -- 
    ra_5261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k2_2067_inst_ack_0, ack => convolve_CP_4643_elements(197)); -- 
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	230 
    -- CP-element group 198: 	244 
    -- CP-element group 198: 	248 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	29 
    -- CP-element group 198: 	195 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k2_2067_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k2_2067_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k2_2067_Update/ca
      -- 
    ca_5266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k2_2067_inst_ack_1, ack => convolve_CP_4643_elements(198)); -- 
    -- CP-element group 199:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	23 
    -- CP-element group 199: marked-predecessors 
    -- CP-element group 199: 	202 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k3_2071_sample_start_
      -- CP-element group 199: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k3_2071_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k3_2071_Sample/rr
      -- 
    rr_5274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(199), ack => RPIPE_xxconvolvexxconv_k3_2071_inst_req_0); -- 
    convolve_cp_element_group_199: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_199"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(23) & convolve_CP_4643_elements(202);
      gj_convolve_cp_element_group_199 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(199), clk => clk, reset => reset); --
    end block;
    -- CP-element group 200:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	26 
    -- CP-element group 200: 	70 
    -- CP-element group 200: 	201 
    -- CP-element group 200: 	51 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	246 
    -- CP-element group 200: 	250 
    -- CP-element group 200: 	238 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: marked-successors 
    -- CP-element group 200: 	66 
    -- CP-element group 200: 	47 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k3_2071_update_start_
      -- CP-element group 200: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k3_2071_Update/$entry
      -- CP-element group 200: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k3_2071_Update/cr
      -- 
    cr_5279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(200), ack => RPIPE_xxconvolvexxconv_k3_2071_inst_req_1); -- 
    convolve_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 1,3 => 15,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(70) & convolve_CP_4643_elements(201) & convolve_CP_4643_elements(51) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250) & convolve_CP_4643_elements(238);
      gj_convolve_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  transition  input  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	200 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k3_2071_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k3_2071_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k3_2071_Sample/ra
      -- 
    ra_5275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k3_2071_inst_ack_0, ack => convolve_CP_4643_elements(201)); -- 
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	200 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	244 
    -- CP-element group 202: 	248 
    -- CP-element group 202: 	237 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	29 
    -- CP-element group 202: 	199 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k3_2071_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k3_2071_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/RPIPE_xxconvolvexxconv_k3_2071_Update/ca
      -- 
    ca_5280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k3_2071_inst_ack_1, ack => convolve_CP_4643_elements(202)); -- 
    -- CP-element group 203:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	70 
    -- CP-element group 203: 	51 
    -- CP-element group 203: marked-predecessors 
    -- CP-element group 203: 	205 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	205 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2075_Sample/req
      -- CP-element group 203: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2075_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2075_Sample/$entry
      -- 
    req_5288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(203), ack => W_read_k_2011_delayed_1_0_2073_inst_req_0); -- 
    convolve_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(70) & convolve_CP_4643_elements(51) & convolve_CP_4643_elements(205);
      gj_convolve_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	26 
    -- CP-element group 204: marked-predecessors 
    -- CP-element group 204: 	224 
    -- CP-element group 204: 	206 
    -- CP-element group 204: 	246 
    -- CP-element group 204: 	250 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	206 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2075_Update/req
      -- CP-element group 204: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2075_Update/$entry
      -- CP-element group 204: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2075_update_start_
      -- 
    req_5293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(204), ack => W_read_k_2011_delayed_1_0_2073_inst_req_1); -- 
    convolve_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(224) & convolve_CP_4643_elements(206) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250);
      gj_convolve_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: successors 
    -- CP-element group 205: marked-successors 
    -- CP-element group 205: 	66 
    -- CP-element group 205: 	47 
    -- CP-element group 205: 	203 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2075_Sample/ack
      -- CP-element group 205: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2075_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2075_Sample/$exit
      -- 
    ack_5289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2011_delayed_1_0_2073_inst_ack_0, ack => convolve_CP_4643_elements(205)); -- 
    -- CP-element group 206:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	204 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	223 
    -- CP-element group 206: 	244 
    -- CP-element group 206: 	248 
    -- CP-element group 206: marked-successors 
    -- CP-element group 206: 	29 
    -- CP-element group 206: 	204 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2075_Update/ack
      -- CP-element group 206: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2075_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2075_update_completed_
      -- 
    ack_5294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2011_delayed_1_0_2073_inst_ack_1, ack => convolve_CP_4643_elements(206)); -- 
    -- CP-element group 207:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	70 
    -- CP-element group 207: 	51 
    -- CP-element group 207: marked-predecessors 
    -- CP-element group 207: 	209 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2084_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2084_Sample/req
      -- CP-element group 207: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2084_sample_start_
      -- 
    req_5302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(207), ack => W_read_k_2017_delayed_1_0_2082_inst_req_0); -- 
    convolve_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(70) & convolve_CP_4643_elements(51) & convolve_CP_4643_elements(209);
      gj_convolve_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	26 
    -- CP-element group 208: marked-predecessors 
    -- CP-element group 208: 	231 
    -- CP-element group 208: 	210 
    -- CP-element group 208: 	246 
    -- CP-element group 208: 	250 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2084_Update/req
      -- CP-element group 208: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2084_update_start_
      -- CP-element group 208: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2084_Update/$entry
      -- 
    req_5307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(208), ack => W_read_k_2017_delayed_1_0_2082_inst_req_1); -- 
    convolve_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(231) & convolve_CP_4643_elements(210) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250);
      gj_convolve_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209: marked-successors 
    -- CP-element group 209: 	66 
    -- CP-element group 209: 	47 
    -- CP-element group 209: 	207 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2084_Sample/$exit
      -- CP-element group 209: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2084_Sample/ack
      -- CP-element group 209: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2084_sample_completed_
      -- 
    ack_5303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2017_delayed_1_0_2082_inst_ack_0, ack => convolve_CP_4643_elements(209)); -- 
    -- CP-element group 210:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	230 
    -- CP-element group 210: 	244 
    -- CP-element group 210: 	248 
    -- CP-element group 210: marked-successors 
    -- CP-element group 210: 	29 
    -- CP-element group 210: 	208 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2084_update_completed_
      -- CP-element group 210: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2084_Update/ack
      -- CP-element group 210: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2084_Update/$exit
      -- 
    ack_5308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2017_delayed_1_0_2082_inst_ack_1, ack => convolve_CP_4643_elements(210)); -- 
    -- CP-element group 211:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	70 
    -- CP-element group 211: 	51 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	213 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2093_sample_start_
      -- CP-element group 211: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2093_Sample/req
      -- CP-element group 211: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2093_Sample/$entry
      -- 
    req_5316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(211), ack => W_read_k_2023_delayed_1_0_2091_inst_req_0); -- 
    convolve_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(70) & convolve_CP_4643_elements(51) & convolve_CP_4643_elements(213);
      gj_convolve_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	26 
    -- CP-element group 212: marked-predecessors 
    -- CP-element group 212: 	214 
    -- CP-element group 212: 	246 
    -- CP-element group 212: 	250 
    -- CP-element group 212: 	238 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	214 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2093_update_start_
      -- CP-element group 212: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2093_Update/req
      -- CP-element group 212: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2093_Update/$entry
      -- 
    req_5321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(212), ack => W_read_k_2023_delayed_1_0_2091_inst_req_1); -- 
    convolve_cp_element_group_212: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_212"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(214) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250) & convolve_CP_4643_elements(238);
      gj_convolve_cp_element_group_212 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(212), clk => clk, reset => reset); --
    end block;
    -- CP-element group 213:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: marked-successors 
    -- CP-element group 213: 	66 
    -- CP-element group 213: 	47 
    -- CP-element group 213: 	211 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2093_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2093_Sample/ack
      -- CP-element group 213: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2093_Sample/$exit
      -- 
    ack_5317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2023_delayed_1_0_2091_inst_ack_0, ack => convolve_CP_4643_elements(213)); -- 
    -- CP-element group 214:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	212 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	244 
    -- CP-element group 214: 	248 
    -- CP-element group 214: 	237 
    -- CP-element group 214: marked-successors 
    -- CP-element group 214: 	29 
    -- CP-element group 214: 	212 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2093_Update/ack
      -- CP-element group 214: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2093_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2093_update_completed_
      -- 
    ack_5322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2023_delayed_1_0_2091_inst_ack_1, ack => convolve_CP_4643_elements(214)); -- 
    -- CP-element group 215:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	32 
    -- CP-element group 215: marked-predecessors 
    -- CP-element group 215: 	217 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	217 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2132_Sample/req
      -- CP-element group 215: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2132_Sample/$entry
      -- CP-element group 215: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2132_sample_start_
      -- 
    req_5330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(215), ack => W_acc_2059_delayed_1_0_2130_inst_req_0); -- 
    convolve_cp_element_group_215: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_215"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(32) & convolve_CP_4643_elements(217);
      gj_convolve_cp_element_group_215 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(215), clk => clk, reset => reset); --
    end block;
    -- CP-element group 216:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	26 
    -- CP-element group 216: marked-predecessors 
    -- CP-element group 216: 	246 
    -- CP-element group 216: 	250 
    -- CP-element group 216: 	218 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	218 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2132_Update/$entry
      -- CP-element group 216: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2132_Update/req
      -- CP-element group 216: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2132_update_start_
      -- 
    req_5335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(216), ack => W_acc_2059_delayed_1_0_2130_inst_req_1); -- 
    convolve_cp_element_group_216: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_216"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(246) & convolve_CP_4643_elements(250) & convolve_CP_4643_elements(218);
      gj_convolve_cp_element_group_216 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(216), clk => clk, reset => reset); --
    end block;
    -- CP-element group 217:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	215 
    -- CP-element group 217: successors 
    -- CP-element group 217: marked-successors 
    -- CP-element group 217: 	30 
    -- CP-element group 217: 	215 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2132_Sample/ack
      -- CP-element group 217: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2132_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2132_sample_completed_
      -- 
    ack_5331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc_2059_delayed_1_0_2130_inst_ack_0, ack => convolve_CP_4643_elements(217)); -- 
    -- CP-element group 218:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	216 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	244 
    -- CP-element group 218: 	248 
    -- CP-element group 218: marked-successors 
    -- CP-element group 218: 	29 
    -- CP-element group 218: 	216 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2132_Update/ack
      -- CP-element group 218: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2132_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2132_update_completed_
      -- 
    ack_5336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc_2059_delayed_1_0_2130_inst_ack_1, ack => convolve_CP_4643_elements(218)); -- 
    -- CP-element group 219:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	70 
    -- CP-element group 219: 	51 
    -- CP-element group 219: marked-predecessors 
    -- CP-element group 219: 	221 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2182_sample_start_
      -- CP-element group 219: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2182_Sample/$entry
      -- CP-element group 219: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2182_Sample/req
      -- 
    req_5344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(219), ack => W_store_kernel_2105_delayed_1_0_2180_inst_req_0); -- 
    convolve_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(70) & convolve_CP_4643_elements(51) & convolve_CP_4643_elements(221);
      gj_convolve_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: marked-predecessors 
    -- CP-element group 220: 	222 
    -- CP-element group 220: 	224 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	222 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2182_Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2182_update_start_
      -- CP-element group 220: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2182_Update/req
      -- 
    req_5349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(220), ack => W_store_kernel_2105_delayed_1_0_2180_inst_req_1); -- 
    convolve_cp_element_group_220: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_220"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(222) & convolve_CP_4643_elements(224);
      gj_convolve_cp_element_group_220 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(220), clk => clk, reset => reset); --
    end block;
    -- CP-element group 221:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: marked-successors 
    -- CP-element group 221: 	66 
    -- CP-element group 221: 	47 
    -- CP-element group 221: 	219 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2182_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2182_Sample/ack
      -- CP-element group 221: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2182_Sample/$exit
      -- 
    ack_5345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2105_delayed_1_0_2180_inst_ack_0, ack => convolve_CP_4643_elements(221)); -- 
    -- CP-element group 222:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	220 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222: marked-successors 
    -- CP-element group 222: 	220 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2182_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2182_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2182_Update/ack
      -- 
    ack_5350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2105_delayed_1_0_2180_inst_ack_1, ack => convolve_CP_4643_elements(222)); -- 
    -- CP-element group 223:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	194 
    -- CP-element group 223: 	222 
    -- CP-element group 223: 	182 
    -- CP-element group 223: 	206 
    -- CP-element group 223: marked-predecessors 
    -- CP-element group 223: 	225 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k1_2184_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k1_2184_Sample/req
      -- CP-element group 223: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k1_2184_Sample/$entry
      -- 
    req_5358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(223), ack => WPIPE_xxconvolvexxconv_k1_2184_inst_req_0); -- 
    convolve_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(194) & convolve_CP_4643_elements(222) & convolve_CP_4643_elements(182) & convolve_CP_4643_elements(206) & convolve_CP_4643_elements(225);
      gj_convolve_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	225 
    -- CP-element group 224: marked-successors 
    -- CP-element group 224: 	192 
    -- CP-element group 224: 	204 
    -- CP-element group 224: 	180 
    -- CP-element group 224: 	220 
    -- CP-element group 224:  members (6) 
      -- CP-element group 224: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k1_2184_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k1_2184_update_start_
      -- CP-element group 224: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k1_2184_Update/req
      -- CP-element group 224: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k1_2184_Update/$entry
      -- CP-element group 224: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k1_2184_Sample/ack
      -- CP-element group 224: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k1_2184_Sample/$exit
      -- 
    ack_5359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k1_2184_inst_ack_0, ack => convolve_CP_4643_elements(224)); -- 
    req_5363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(224), ack => WPIPE_xxconvolvexxconv_k1_2184_inst_req_1); -- 
    -- CP-element group 225:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	224 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	275 
    -- CP-element group 225: marked-successors 
    -- CP-element group 225: 	223 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k1_2184_Update/ack
      -- CP-element group 225: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k1_2184_Update/$exit
      -- CP-element group 225: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k1_2184_update_completed_
      -- 
    ack_5364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k1_2184_inst_ack_1, ack => convolve_CP_4643_elements(225)); -- 
    -- CP-element group 226:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	70 
    -- CP-element group 226: 	51 
    -- CP-element group 226: marked-predecessors 
    -- CP-element group 226: 	228 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	228 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2189_Sample/req
      -- CP-element group 226: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2189_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2189_sample_start_
      -- 
    req_5372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(226), ack => W_store_kernel_2109_delayed_1_0_2187_inst_req_0); -- 
    convolve_cp_element_group_226: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_226"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(70) & convolve_CP_4643_elements(51) & convolve_CP_4643_elements(228);
      gj_convolve_cp_element_group_226 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 227:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: marked-predecessors 
    -- CP-element group 227: 	229 
    -- CP-element group 227: 	231 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	229 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2189_Update/req
      -- CP-element group 227: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2189_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2189_update_start_
      -- 
    req_5377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(227), ack => W_store_kernel_2109_delayed_1_0_2187_inst_req_1); -- 
    convolve_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(229) & convolve_CP_4643_elements(231);
      gj_convolve_cp_element_group_227 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: successors 
    -- CP-element group 228: marked-successors 
    -- CP-element group 228: 	66 
    -- CP-element group 228: 	226 
    -- CP-element group 228: 	47 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2189_Sample/ack
      -- CP-element group 228: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2189_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2189_sample_completed_
      -- 
    ack_5373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2109_delayed_1_0_2187_inst_ack_0, ack => convolve_CP_4643_elements(228)); -- 
    -- CP-element group 229:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229: marked-successors 
    -- CP-element group 229: 	227 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2189_Update/ack
      -- CP-element group 229: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2189_Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2189_update_completed_
      -- 
    ack_5378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2109_delayed_1_0_2187_inst_ack_1, ack => convolve_CP_4643_elements(229)); -- 
    -- CP-element group 230:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	198 
    -- CP-element group 230: 	229 
    -- CP-element group 230: 	186 
    -- CP-element group 230: 	210 
    -- CP-element group 230: marked-predecessors 
    -- CP-element group 230: 	232 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k2_2191_Sample/req
      -- CP-element group 230: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k2_2191_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k2_2191_sample_start_
      -- 
    req_5386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(230), ack => WPIPE_xxconvolvexxconv_k2_2191_inst_req_0); -- 
    convolve_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(198) & convolve_CP_4643_elements(229) & convolve_CP_4643_elements(186) & convolve_CP_4643_elements(210) & convolve_CP_4643_elements(232);
      gj_convolve_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231: marked-successors 
    -- CP-element group 231: 	196 
    -- CP-element group 231: 	227 
    -- CP-element group 231: 	184 
    -- CP-element group 231: 	208 
    -- CP-element group 231:  members (6) 
      -- CP-element group 231: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k2_2191_Update/req
      -- CP-element group 231: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k2_2191_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k2_2191_Sample/ack
      -- CP-element group 231: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k2_2191_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k2_2191_update_start_
      -- CP-element group 231: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k2_2191_sample_completed_
      -- 
    ack_5387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k2_2191_inst_ack_0, ack => convolve_CP_4643_elements(231)); -- 
    req_5391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(231), ack => WPIPE_xxconvolvexxconv_k2_2191_inst_req_1); -- 
    -- CP-element group 232:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	275 
    -- CP-element group 232: marked-successors 
    -- CP-element group 232: 	230 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k2_2191_Update/ack
      -- CP-element group 232: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k2_2191_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k2_2191_update_completed_
      -- 
    ack_5392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k2_2191_inst_ack_1, ack => convolve_CP_4643_elements(232)); -- 
    -- CP-element group 233:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	70 
    -- CP-element group 233: 	51 
    -- CP-element group 233: marked-predecessors 
    -- CP-element group 233: 	235 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2196_Sample/$entry
      -- CP-element group 233: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2196_Sample/req
      -- CP-element group 233: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2196_sample_start_
      -- 
    req_5400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(233), ack => W_store_kernel_2113_delayed_1_0_2194_inst_req_0); -- 
    convolve_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(70) & convolve_CP_4643_elements(51) & convolve_CP_4643_elements(235);
      gj_convolve_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: marked-predecessors 
    -- CP-element group 234: 	236 
    -- CP-element group 234: 	238 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2196_Update/req
      -- CP-element group 234: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2196_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2196_update_start_
      -- 
    req_5405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(234), ack => W_store_kernel_2113_delayed_1_0_2194_inst_req_1); -- 
    convolve_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(236) & convolve_CP_4643_elements(238);
      gj_convolve_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: marked-successors 
    -- CP-element group 235: 	66 
    -- CP-element group 235: 	47 
    -- CP-element group 235: 	233 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2196_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2196_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2196_sample_completed_
      -- 
    ack_5401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2113_delayed_1_0_2194_inst_ack_0, ack => convolve_CP_4643_elements(235)); -- 
    -- CP-element group 236:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236: marked-successors 
    -- CP-element group 236: 	234 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2196_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2196_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2196_Update/ack
      -- 
    ack_5406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2113_delayed_1_0_2194_inst_ack_1, ack => convolve_CP_4643_elements(236)); -- 
    -- CP-element group 237:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	190 
    -- CP-element group 237: 	202 
    -- CP-element group 237: 	214 
    -- CP-element group 237: 	236 
    -- CP-element group 237: marked-predecessors 
    -- CP-element group 237: 	239 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k3_2198_Sample/req
      -- CP-element group 237: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k3_2198_Sample/$entry
      -- CP-element group 237: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k3_2198_sample_start_
      -- 
    req_5414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(237), ack => WPIPE_xxconvolvexxconv_k3_2198_inst_req_0); -- 
    convolve_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(190) & convolve_CP_4643_elements(202) & convolve_CP_4643_elements(214) & convolve_CP_4643_elements(236) & convolve_CP_4643_elements(239);
      gj_convolve_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238: marked-successors 
    -- CP-element group 238: 	200 
    -- CP-element group 238: 	188 
    -- CP-element group 238: 	212 
    -- CP-element group 238: 	234 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k3_2198_sample_completed_
      -- CP-element group 238: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k3_2198_update_start_
      -- CP-element group 238: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k3_2198_Sample/ack
      -- CP-element group 238: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k3_2198_Sample/$exit
      -- CP-element group 238: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k3_2198_Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k3_2198_Update/req
      -- 
    ack_5415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k3_2198_inst_ack_0, ack => convolve_CP_4643_elements(238)); -- 
    req_5419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(238), ack => WPIPE_xxconvolvexxconv_k3_2198_inst_req_1); -- 
    -- CP-element group 239:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	275 
    -- CP-element group 239: marked-successors 
    -- CP-element group 239: 	237 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k3_2198_update_completed_
      -- CP-element group 239: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k3_2198_Update/$exit
      -- CP-element group 239: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_xxconvolvexxconv_k3_2198_Update/ack
      -- 
    ack_5420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k3_2198_inst_ack_1, ack => convolve_CP_4643_elements(239)); -- 
    -- CP-element group 240:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	89 
    -- CP-element group 240: 	108 
    -- CP-element group 240: marked-predecessors 
    -- CP-element group 240: 	242 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	242 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2241_Sample/req
      -- CP-element group 240: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2241_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2241_sample_start_
      -- 
    req_5428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(240), ack => W_num_done_2156_delayed_1_0_2239_inst_req_0); -- 
    convolve_cp_element_group_240: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_240"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(89) & convolve_CP_4643_elements(108) & convolve_CP_4643_elements(242);
      gj_convolve_cp_element_group_240 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(240), clk => clk, reset => reset); --
    end block;
    -- CP-element group 241:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	26 
    -- CP-element group 241: marked-predecessors 
    -- CP-element group 241: 	243 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2241_Update/req
      -- CP-element group 241: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2241_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2241_update_start_
      -- 
    req_5433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(241), ack => W_num_done_2156_delayed_1_0_2239_inst_req_1); -- 
    convolve_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(243);
      gj_convolve_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	240 
    -- CP-element group 242: successors 
    -- CP-element group 242: marked-successors 
    -- CP-element group 242: 	85 
    -- CP-element group 242: 	104 
    -- CP-element group 242: 	240 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2241_Sample/ack
      -- CP-element group 242: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2241_Sample/$exit
      -- CP-element group 242: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2241_sample_completed_
      -- 
    ack_5429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2156_delayed_1_0_2239_inst_ack_0, ack => convolve_CP_4643_elements(242)); -- 
    -- CP-element group 243:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	275 
    -- CP-element group 243: marked-successors 
    -- CP-element group 243: 	29 
    -- CP-element group 243: 	241 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2241_Update/ack
      -- CP-element group 243: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2241_Update/$exit
      -- CP-element group 243: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2241_update_completed_
      -- 
    ack_5434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2156_delayed_1_0_2239_inst_ack_1, ack => convolve_CP_4643_elements(243)); -- 
    -- CP-element group 244:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	125 
    -- CP-element group 244: 	129 
    -- CP-element group 244: 	133 
    -- CP-element group 244: 	137 
    -- CP-element group 244: 	141 
    -- CP-element group 244: 	190 
    -- CP-element group 244: 	194 
    -- CP-element group 244: 	198 
    -- CP-element group 244: 	145 
    -- CP-element group 244: 	149 
    -- CP-element group 244: 	153 
    -- CP-element group 244: 	157 
    -- CP-element group 244: 	182 
    -- CP-element group 244: 	186 
    -- CP-element group 244: 	202 
    -- CP-element group 244: 	206 
    -- CP-element group 244: 	210 
    -- CP-element group 244: 	214 
    -- CP-element group 244: 	218 
    -- CP-element group 244: marked-predecessors 
    -- CP-element group 244: 	246 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	246 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2250_Sample/rr
      -- CP-element group 244: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2250_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2250_sample_start_
      -- 
    rr_5442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(244), ack => slice_2250_inst_req_0); -- 
    convolve_cp_element_group_244: block -- 
      constant place_capacities: IntegerArray(0 to 19) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1);
      constant place_markings: IntegerArray(0 to 19)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 1);
      constant place_delays: IntegerArray(0 to 19) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_244"; 
      signal preds: BooleanArray(1 to 20); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(125) & convolve_CP_4643_elements(129) & convolve_CP_4643_elements(133) & convolve_CP_4643_elements(137) & convolve_CP_4643_elements(141) & convolve_CP_4643_elements(190) & convolve_CP_4643_elements(194) & convolve_CP_4643_elements(198) & convolve_CP_4643_elements(145) & convolve_CP_4643_elements(149) & convolve_CP_4643_elements(153) & convolve_CP_4643_elements(157) & convolve_CP_4643_elements(182) & convolve_CP_4643_elements(186) & convolve_CP_4643_elements(202) & convolve_CP_4643_elements(206) & convolve_CP_4643_elements(210) & convolve_CP_4643_elements(214) & convolve_CP_4643_elements(218) & convolve_CP_4643_elements(246);
      gj_convolve_cp_element_group_244 : generic_join generic map(name => joinName, number_of_predecessors => 20, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(244), clk => clk, reset => reset); --
    end block;
    -- CP-element group 245:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: marked-predecessors 
    -- CP-element group 245: 	247 
    -- CP-element group 245: 	258 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2250_Update/cr
      -- CP-element group 245: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2250_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2250_update_start_
      -- 
    cr_5447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(245), ack => slice_2250_inst_req_1); -- 
    convolve_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(247) & convolve_CP_4643_elements(258);
      gj_convolve_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	244 
    -- CP-element group 246: successors 
    -- CP-element group 246: marked-successors 
    -- CP-element group 246: 	123 
    -- CP-element group 246: 	127 
    -- CP-element group 246: 	131 
    -- CP-element group 246: 	135 
    -- CP-element group 246: 	139 
    -- CP-element group 246: 	143 
    -- CP-element group 246: 	192 
    -- CP-element group 246: 	196 
    -- CP-element group 246: 	200 
    -- CP-element group 246: 	147 
    -- CP-element group 246: 	151 
    -- CP-element group 246: 	155 
    -- CP-element group 246: 	184 
    -- CP-element group 246: 	188 
    -- CP-element group 246: 	204 
    -- CP-element group 246: 	208 
    -- CP-element group 246: 	212 
    -- CP-element group 246: 	180 
    -- CP-element group 246: 	244 
    -- CP-element group 246: 	216 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2250_Sample/ra
      -- CP-element group 246: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2250_Sample/$exit
      -- CP-element group 246: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2250_sample_completed_
      -- 
    ra_5443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2250_inst_ack_0, ack => convolve_CP_4643_elements(246)); -- 
    -- CP-element group 247:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	256 
    -- CP-element group 247: marked-successors 
    -- CP-element group 247: 	245 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2250_Update/ca
      -- CP-element group 247: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2250_Update/$exit
      -- CP-element group 247: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2250_update_completed_
      -- 
    ca_5448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2250_inst_ack_1, ack => convolve_CP_4643_elements(247)); -- 
    -- CP-element group 248:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	125 
    -- CP-element group 248: 	129 
    -- CP-element group 248: 	133 
    -- CP-element group 248: 	137 
    -- CP-element group 248: 	141 
    -- CP-element group 248: 	190 
    -- CP-element group 248: 	194 
    -- CP-element group 248: 	198 
    -- CP-element group 248: 	145 
    -- CP-element group 248: 	149 
    -- CP-element group 248: 	153 
    -- CP-element group 248: 	157 
    -- CP-element group 248: 	182 
    -- CP-element group 248: 	186 
    -- CP-element group 248: 	202 
    -- CP-element group 248: 	206 
    -- CP-element group 248: 	210 
    -- CP-element group 248: 	214 
    -- CP-element group 248: 	218 
    -- CP-element group 248: marked-predecessors 
    -- CP-element group 248: 	250 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	250 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2254_Sample/rr
      -- CP-element group 248: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2254_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2254_sample_start_
      -- 
    rr_5456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(248), ack => slice_2254_inst_req_0); -- 
    convolve_cp_element_group_248: block -- 
      constant place_capacities: IntegerArray(0 to 19) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1);
      constant place_markings: IntegerArray(0 to 19)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 1);
      constant place_delays: IntegerArray(0 to 19) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_248"; 
      signal preds: BooleanArray(1 to 20); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(125) & convolve_CP_4643_elements(129) & convolve_CP_4643_elements(133) & convolve_CP_4643_elements(137) & convolve_CP_4643_elements(141) & convolve_CP_4643_elements(190) & convolve_CP_4643_elements(194) & convolve_CP_4643_elements(198) & convolve_CP_4643_elements(145) & convolve_CP_4643_elements(149) & convolve_CP_4643_elements(153) & convolve_CP_4643_elements(157) & convolve_CP_4643_elements(182) & convolve_CP_4643_elements(186) & convolve_CP_4643_elements(202) & convolve_CP_4643_elements(206) & convolve_CP_4643_elements(210) & convolve_CP_4643_elements(214) & convolve_CP_4643_elements(218) & convolve_CP_4643_elements(250);
      gj_convolve_cp_element_group_248 : generic_join generic map(name => joinName, number_of_predecessors => 20, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(248), clk => clk, reset => reset); --
    end block;
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	251 
    -- CP-element group 249: 	269 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2254_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2254_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2254_update_start_
      -- 
    cr_5461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(249), ack => slice_2254_inst_req_1); -- 
    convolve_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(251) & convolve_CP_4643_elements(269);
      gj_convolve_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	248 
    -- CP-element group 250: successors 
    -- CP-element group 250: marked-successors 
    -- CP-element group 250: 	123 
    -- CP-element group 250: 	127 
    -- CP-element group 250: 	131 
    -- CP-element group 250: 	135 
    -- CP-element group 250: 	139 
    -- CP-element group 250: 	143 
    -- CP-element group 250: 	192 
    -- CP-element group 250: 	196 
    -- CP-element group 250: 	200 
    -- CP-element group 250: 	147 
    -- CP-element group 250: 	151 
    -- CP-element group 250: 	155 
    -- CP-element group 250: 	184 
    -- CP-element group 250: 	188 
    -- CP-element group 250: 	204 
    -- CP-element group 250: 	208 
    -- CP-element group 250: 	212 
    -- CP-element group 250: 	180 
    -- CP-element group 250: 	248 
    -- CP-element group 250: 	216 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2254_Sample/ra
      -- CP-element group 250: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2254_Sample/$exit
      -- CP-element group 250: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2254_sample_completed_
      -- 
    ra_5457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2254_inst_ack_0, ack => convolve_CP_4643_elements(250)); -- 
    -- CP-element group 251:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	267 
    -- CP-element group 251: marked-successors 
    -- CP-element group 251: 	249 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2254_Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2254_Update/ca
      -- CP-element group 251: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/slice_2254_update_completed_
      -- 
    ca_5462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2254_inst_ack_1, ack => convolve_CP_4643_elements(251)); -- 
    -- CP-element group 252:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	89 
    -- CP-element group 252: 	108 
    -- CP-element group 252: marked-predecessors 
    -- CP-element group 252: 	254 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	254 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2258_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2258_Sample/req
      -- CP-element group 252: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2258_Sample/$entry
      -- 
    req_5470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(252), ack => W_num_done_2169_delayed_2_0_2256_inst_req_0); -- 
    convolve_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(89) & convolve_CP_4643_elements(108) & convolve_CP_4643_elements(254);
      gj_convolve_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: marked-predecessors 
    -- CP-element group 253: 	255 
    -- CP-element group 253: 	258 
    -- CP-element group 253: 	261 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2258_update_start_
      -- CP-element group 253: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2258_Update/req
      -- CP-element group 253: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2258_Update/$entry
      -- 
    req_5475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(253), ack => W_num_done_2169_delayed_2_0_2256_inst_req_1); -- 
    convolve_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(255) & convolve_CP_4643_elements(258) & convolve_CP_4643_elements(261);
      gj_convolve_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	252 
    -- CP-element group 254: successors 
    -- CP-element group 254: marked-successors 
    -- CP-element group 254: 	85 
    -- CP-element group 254: 	104 
    -- CP-element group 254: 	252 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2258_sample_completed_
      -- CP-element group 254: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2258_Sample/ack
      -- CP-element group 254: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2258_Sample/$exit
      -- 
    ack_5471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2169_delayed_2_0_2256_inst_ack_0, ack => convolve_CP_4643_elements(254)); -- 
    -- CP-element group 255:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255: 	260 
    -- CP-element group 255: marked-successors 
    -- CP-element group 255: 	253 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2258_update_completed_
      -- CP-element group 255: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2258_Update/ack
      -- CP-element group 255: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2258_Update/$exit
      -- 
    ack_5476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2169_delayed_2_0_2256_inst_ack_1, ack => convolve_CP_4643_elements(255)); -- 
    -- CP-element group 256:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	247 
    -- CP-element group 256: 	255 
    -- CP-element group 256: marked-predecessors 
    -- CP-element group 256: 	258 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	258 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2262_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2262_Sample/rr
      -- CP-element group 256: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2262_Sample/$entry
      -- 
    rr_5484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(256), ack => type_cast_2262_inst_req_0); -- 
    convolve_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(247) & convolve_CP_4643_elements(255) & convolve_CP_4643_elements(258);
      gj_convolve_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: marked-predecessors 
    -- CP-element group 257: 	259 
    -- CP-element group 257: 	261 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2262_update_start_
      -- CP-element group 257: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2262_Update/cr
      -- CP-element group 257: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2262_Update/$entry
      -- 
    cr_5489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(257), ack => type_cast_2262_inst_req_1); -- 
    convolve_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(259) & convolve_CP_4643_elements(261);
      gj_convolve_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	256 
    -- CP-element group 258: successors 
    -- CP-element group 258: marked-successors 
    -- CP-element group 258: 	245 
    -- CP-element group 258: 	253 
    -- CP-element group 258: 	256 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2262_sample_completed_
      -- CP-element group 258: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2262_Sample/ra
      -- CP-element group 258: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2262_Sample/$exit
      -- 
    ra_5485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2262_inst_ack_0, ack => convolve_CP_4643_elements(258)); -- 
    -- CP-element group 259:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	257 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2262_update_completed_
      -- CP-element group 259: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2262_Update/ca
      -- CP-element group 259: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2262_Update/$exit
      -- 
    ca_5490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2262_inst_ack_1, ack => convolve_CP_4643_elements(259)); -- 
    -- CP-element group 260:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	255 
    -- CP-element group 260: 	259 
    -- CP-element group 260: marked-predecessors 
    -- CP-element group 260: 	273 
    -- CP-element group 260: 	262 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2260_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2260_Sample/req
      -- CP-element group 260: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2260_Sample/$entry
      -- 
    req_5498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(260), ack => WPIPE_maxpool_output_pipe_2260_inst_req_0); -- 
    convolve_cp_element_group_260: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_260"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(255) & convolve_CP_4643_elements(259) & convolve_CP_4643_elements(273) & convolve_CP_4643_elements(262);
      gj_convolve_cp_element_group_260 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(260), clk => clk, reset => reset); --
    end block;
    -- CP-element group 261:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261: marked-successors 
    -- CP-element group 261: 	253 
    -- CP-element group 261: 	257 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2260_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2260_sample_completed_
      -- CP-element group 261: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2260_Sample/ack
      -- CP-element group 261: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2260_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2260_Update/req
      -- CP-element group 261: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2260_update_start_
      -- 
    ack_5499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2260_inst_ack_0, ack => convolve_CP_4643_elements(261)); -- 
    req_5503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(261), ack => WPIPE_maxpool_output_pipe_2260_inst_req_1); -- 
    -- CP-element group 262:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	271 
    -- CP-element group 262: marked-successors 
    -- CP-element group 262: 	260 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2260_Update/ack
      -- CP-element group 262: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2260_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2260_update_completed_
      -- 
    ack_5504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2260_inst_ack_1, ack => convolve_CP_4643_elements(262)); -- 
    -- CP-element group 263:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	89 
    -- CP-element group 263: 	108 
    -- CP-element group 263: marked-predecessors 
    -- CP-element group 263: 	265 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	265 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2266_sample_start_
      -- CP-element group 263: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2266_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2266_Sample/req
      -- 
    req_5512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(263), ack => W_num_done_2174_delayed_2_0_2264_inst_req_0); -- 
    convolve_cp_element_group_263: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_263"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(89) & convolve_CP_4643_elements(108) & convolve_CP_4643_elements(265);
      gj_convolve_cp_element_group_263 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(263), clk => clk, reset => reset); --
    end block;
    -- CP-element group 264:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: marked-predecessors 
    -- CP-element group 264: 	266 
    -- CP-element group 264: 	269 
    -- CP-element group 264: 	272 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	266 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2266_Update/req
      -- CP-element group 264: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2266_Update/$entry
      -- CP-element group 264: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2266_update_start_
      -- 
    req_5517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(264), ack => W_num_done_2174_delayed_2_0_2264_inst_req_1); -- 
    convolve_cp_element_group_264: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_264"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(266) & convolve_CP_4643_elements(269) & convolve_CP_4643_elements(272);
      gj_convolve_cp_element_group_264 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(264), clk => clk, reset => reset); --
    end block;
    -- CP-element group 265:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	263 
    -- CP-element group 265: successors 
    -- CP-element group 265: marked-successors 
    -- CP-element group 265: 	85 
    -- CP-element group 265: 	104 
    -- CP-element group 265: 	263 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2266_sample_completed_
      -- CP-element group 265: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2266_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2266_Sample/ack
      -- 
    ack_5513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2174_delayed_2_0_2264_inst_ack_0, ack => convolve_CP_4643_elements(265)); -- 
    -- CP-element group 266:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	264 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266: 	271 
    -- CP-element group 266: marked-successors 
    -- CP-element group 266: 	264 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2266_Update/ack
      -- CP-element group 266: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2266_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/assign_stmt_2266_update_completed_
      -- 
    ack_5518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2174_delayed_2_0_2264_inst_ack_1, ack => convolve_CP_4643_elements(266)); -- 
    -- CP-element group 267:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	251 
    -- CP-element group 267: 	266 
    -- CP-element group 267: marked-predecessors 
    -- CP-element group 267: 	269 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	269 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2270_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2270_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2270_Sample/rr
      -- 
    rr_5526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(267), ack => type_cast_2270_inst_req_0); -- 
    convolve_cp_element_group_267: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_267"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(251) & convolve_CP_4643_elements(266) & convolve_CP_4643_elements(269);
      gj_convolve_cp_element_group_267 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(267), clk => clk, reset => reset); --
    end block;
    -- CP-element group 268:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: marked-predecessors 
    -- CP-element group 268: 	270 
    -- CP-element group 268: 	272 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	270 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2270_update_start_
      -- CP-element group 268: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2270_Update/$entry
      -- CP-element group 268: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2270_Update/cr
      -- 
    cr_5531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(268), ack => type_cast_2270_inst_req_1); -- 
    convolve_cp_element_group_268: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_268"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(270) & convolve_CP_4643_elements(272);
      gj_convolve_cp_element_group_268 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(268), clk => clk, reset => reset); --
    end block;
    -- CP-element group 269:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	267 
    -- CP-element group 269: successors 
    -- CP-element group 269: marked-successors 
    -- CP-element group 269: 	249 
    -- CP-element group 269: 	267 
    -- CP-element group 269: 	264 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2270_Sample/ra
      -- CP-element group 269: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2270_sample_completed_
      -- CP-element group 269: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2270_Sample/$exit
      -- 
    ra_5527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2270_inst_ack_0, ack => convolve_CP_4643_elements(269)); -- 
    -- CP-element group 270:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	268 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270: marked-successors 
    -- CP-element group 270: 	268 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2270_update_completed_
      -- CP-element group 270: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2270_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/type_cast_2270_Update/ca
      -- 
    ca_5532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2270_inst_ack_1, ack => convolve_CP_4643_elements(270)); -- 
    -- CP-element group 271:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	266 
    -- CP-element group 271: 	270 
    -- CP-element group 271: 	262 
    -- CP-element group 271: marked-predecessors 
    -- CP-element group 271: 	273 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2268_sample_start_
      -- CP-element group 271: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2268_Sample/$entry
      -- CP-element group 271: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2268_Sample/req
      -- 
    req_5540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(271), ack => WPIPE_maxpool_output_pipe_2268_inst_req_0); -- 
    convolve_cp_element_group_271: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_271"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(266) & convolve_CP_4643_elements(270) & convolve_CP_4643_elements(262) & convolve_CP_4643_elements(273);
      gj_convolve_cp_element_group_271 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(271), clk => clk, reset => reset); --
    end block;
    -- CP-element group 272:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272: marked-successors 
    -- CP-element group 272: 	268 
    -- CP-element group 272: 	264 
    -- CP-element group 272:  members (6) 
      -- CP-element group 272: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2268_Sample/ack
      -- CP-element group 272: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2268_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2268_Update/req
      -- CP-element group 272: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2268_sample_completed_
      -- CP-element group 272: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2268_update_start_
      -- CP-element group 272: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2268_Sample/$exit
      -- 
    ack_5541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2268_inst_ack_0, ack => convolve_CP_4643_elements(272)); -- 
    req_5545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(272), ack => WPIPE_maxpool_output_pipe_2268_inst_req_1); -- 
    -- CP-element group 273:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273: marked-successors 
    -- CP-element group 273: 	271 
    -- CP-element group 273: 	260 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2268_Update/$exit
      -- CP-element group 273: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2268_Update/ack
      -- CP-element group 273: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/WPIPE_maxpool_output_pipe_2268_update_completed_
      -- 
    ack_5546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_2268_inst_ack_1, ack => convolve_CP_4643_elements(273)); -- 
    -- CP-element group 274:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	23 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	24 
    -- CP-element group 274:  members (1) 
      -- CP-element group 274: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group convolve_CP_4643_elements(274) is a control-delay.
    cp_element_274_delay: control_delay_element  generic map(name => " 274_delay", delay_value => 1)  port map(req => convolve_CP_4643_elements(23), ack => convolve_CP_4643_elements(274), clk => clk, reset =>reset);
    -- CP-element group 275:  join  transition  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	26 
    -- CP-element group 275: 	225 
    -- CP-element group 275: 	164 
    -- CP-element group 275: 	171 
    -- CP-element group 275: 	232 
    -- CP-element group 275: 	178 
    -- CP-element group 275: 	239 
    -- CP-element group 275: 	243 
    -- CP-element group 275: 	273 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	20 
    -- CP-element group 275:  members (1) 
      -- CP-element group 275: 	 branch_block_stmt_1891/do_while_stmt_1908/do_while_stmt_1908_loop_body/$exit
      -- 
    convolve_cp_element_group_275: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_275"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolve_CP_4643_elements(26) & convolve_CP_4643_elements(225) & convolve_CP_4643_elements(164) & convolve_CP_4643_elements(171) & convolve_CP_4643_elements(232) & convolve_CP_4643_elements(178) & convolve_CP_4643_elements(239) & convolve_CP_4643_elements(243) & convolve_CP_4643_elements(273);
      gj_convolve_cp_element_group_275 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4643_elements(275), clk => clk, reset => reset); --
    end block;
    -- CP-element group 276:  transition  input  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	19 
    -- CP-element group 276: successors 
    -- CP-element group 276:  members (2) 
      -- CP-element group 276: 	 branch_block_stmt_1891/do_while_stmt_1908/loop_exit/$exit
      -- CP-element group 276: 	 branch_block_stmt_1891/do_while_stmt_1908/loop_exit/ack
      -- 
    ack_5551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1908_branch_ack_0, ack => convolve_CP_4643_elements(276)); -- 
    -- CP-element group 277:  transition  input  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	19 
    -- CP-element group 277: successors 
    -- CP-element group 277:  members (2) 
      -- CP-element group 277: 	 branch_block_stmt_1891/do_while_stmt_1908/loop_taken/$exit
      -- CP-element group 277: 	 branch_block_stmt_1891/do_while_stmt_1908/loop_taken/ack
      -- 
    ack_5555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1908_branch_ack_1, ack => convolve_CP_4643_elements(277)); -- 
    -- CP-element group 278:  transition  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	17 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	2 
    -- CP-element group 278:  members (1) 
      -- CP-element group 278: 	 branch_block_stmt_1891/do_while_stmt_1908/$exit
      -- 
    convolve_CP_4643_elements(278) <= convolve_CP_4643_elements(17);
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	2 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_1891/assign_stmt_2277/WPIPE_input_done_pipe_2275_sample_completed_
      -- CP-element group 279: 	 branch_block_stmt_1891/assign_stmt_2277/WPIPE_input_done_pipe_2275_update_start_
      -- CP-element group 279: 	 branch_block_stmt_1891/assign_stmt_2277/WPIPE_input_done_pipe_2275_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_1891/assign_stmt_2277/WPIPE_input_done_pipe_2275_Sample/ack
      -- CP-element group 279: 	 branch_block_stmt_1891/assign_stmt_2277/WPIPE_input_done_pipe_2275_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_1891/assign_stmt_2277/WPIPE_input_done_pipe_2275_Update/req
      -- 
    ack_5568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_2275_inst_ack_0, ack => convolve_CP_4643_elements(279)); -- 
    req_5572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(279), ack => WPIPE_input_done_pipe_2275_inst_req_1); -- 
    -- CP-element group 280:  transition  place  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (8) 
      -- CP-element group 280: 	 branch_block_stmt_1891/assign_stmt_2277__exit__
      -- CP-element group 280: 	 branch_block_stmt_1891/loopback
      -- CP-element group 280: 	 branch_block_stmt_1891/assign_stmt_2277/$exit
      -- CP-element group 280: 	 branch_block_stmt_1891/assign_stmt_2277/WPIPE_input_done_pipe_2275_update_completed_
      -- CP-element group 280: 	 branch_block_stmt_1891/assign_stmt_2277/WPIPE_input_done_pipe_2275_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_1891/assign_stmt_2277/WPIPE_input_done_pipe_2275_Update/ack
      -- CP-element group 280: 	 branch_block_stmt_1891/loopback_PhiReq/$entry
      -- CP-element group 280: 	 branch_block_stmt_1891/loopback_PhiReq/$exit
      -- 
    ack_5573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_2275_inst_ack_1, ack => convolve_CP_4643_elements(280)); -- 
    -- CP-element group 281:  merge  fork  transition  place  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	0 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	3 
    -- CP-element group 281: 	6 
    -- CP-element group 281: 	10 
    -- CP-element group 281: 	11 
    -- CP-element group 281: 	14 
    -- CP-element group 281:  members (22) 
      -- CP-element group 281: 	 branch_block_stmt_1891/merge_stmt_1892__exit__
      -- CP-element group 281: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907__entry__
      -- CP-element group 281: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/$entry
      -- CP-element group 281: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1896_update_start_
      -- CP-element group 281: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1894_sample_start_
      -- CP-element group 281: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1894_Sample/$entry
      -- CP-element group 281: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_num_out_pipe_1894_Sample/rr
      -- CP-element group 281: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1896_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1896_Update/cr
      -- CP-element group 281: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1901_update_start_
      -- CP-element group 281: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1901_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1901_Update/cr
      -- CP-element group 281: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1906_update_start_
      -- CP-element group 281: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_size_pipe_1904_sample_start_
      -- CP-element group 281: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_size_pipe_1904_Sample/$entry
      -- CP-element group 281: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/RPIPE_size_pipe_1904_Sample/rr
      -- CP-element group 281: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1906_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_1891/assign_stmt_1897_to_assign_stmt_1907/SUB_u16_u16_1906_Update/cr
      -- CP-element group 281: 	 branch_block_stmt_1891/merge_stmt_1892_PhiReqMerge
      -- CP-element group 281: 	 branch_block_stmt_1891/merge_stmt_1892_PhiAck/$entry
      -- CP-element group 281: 	 branch_block_stmt_1891/merge_stmt_1892_PhiAck/$exit
      -- CP-element group 281: 	 branch_block_stmt_1891/merge_stmt_1892_PhiAck/dummy
      -- 
    rr_4674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(281), ack => RPIPE_num_out_pipe_1894_inst_req_0); -- 
    cr_4689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(281), ack => SUB_u16_u16_1896_inst_req_1); -- 
    cr_4717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(281), ack => SUB_u16_u16_1901_inst_req_1); -- 
    rr_4730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(281), ack => RPIPE_size_pipe_1904_inst_req_0); -- 
    cr_4745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4643_elements(281), ack => SUB_u16_u16_1906_inst_req_1); -- 
    convolve_CP_4643_elements(281) <= OrReduce(convolve_CP_4643_elements(0) & convolve_CP_4643_elements(280));
    convolve_do_while_stmt_1908_terminator_5556: loop_terminator -- 
      generic map (name => " convolve_do_while_stmt_1908_terminator_5556", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convolve_CP_4643_elements(20),loop_continue => convolve_CP_4643_elements(277),loop_terminate => convolve_CP_4643_elements(276),loop_back => convolve_CP_4643_elements(18),loop_exit => convolve_CP_4643_elements(17),clk => clk, reset => reset); -- 
    phi_stmt_1910_phi_seq_4810_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4643_elements(35);
      convolve_CP_4643_elements(38)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4643_elements(38);
      convolve_CP_4643_elements(39)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4643_elements(40);
      convolve_CP_4643_elements(36) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4643_elements(33);
      convolve_CP_4643_elements(42)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4643_elements(44);
      convolve_CP_4643_elements(43)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4643_elements(45);
      convolve_CP_4643_elements(34) <= phi_mux_reqs(1);
      phi_stmt_1910_phi_seq_4810 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1910_phi_seq_4810") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4643_elements(25), 
          phi_sample_ack => convolve_CP_4643_elements(31), 
          phi_update_req => convolve_CP_4643_elements(27), 
          phi_update_ack => convolve_CP_4643_elements(32), 
          phi_mux_ack => convolve_CP_4643_elements(37), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1916_phi_seq_4854_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4643_elements(54);
      convolve_CP_4643_elements(57)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4643_elements(57);
      convolve_CP_4643_elements(58)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4643_elements(59);
      convolve_CP_4643_elements(55) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4643_elements(52);
      convolve_CP_4643_elements(61)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4643_elements(63);
      convolve_CP_4643_elements(62)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4643_elements(64);
      convolve_CP_4643_elements(53) <= phi_mux_reqs(1);
      phi_stmt_1916_phi_seq_4854 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1916_phi_seq_4854") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4643_elements(48), 
          phi_sample_ack => convolve_CP_4643_elements(49), 
          phi_update_req => convolve_CP_4643_elements(50), 
          phi_update_ack => convolve_CP_4643_elements(51), 
          phi_mux_ack => convolve_CP_4643_elements(56), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1921_phi_seq_4898_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4643_elements(73);
      convolve_CP_4643_elements(76)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4643_elements(76);
      convolve_CP_4643_elements(77)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4643_elements(78);
      convolve_CP_4643_elements(74) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4643_elements(71);
      convolve_CP_4643_elements(80)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4643_elements(82);
      convolve_CP_4643_elements(81)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4643_elements(83);
      convolve_CP_4643_elements(72) <= phi_mux_reqs(1);
      phi_stmt_1921_phi_seq_4898 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1921_phi_seq_4898") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4643_elements(67), 
          phi_sample_ack => convolve_CP_4643_elements(68), 
          phi_update_req => convolve_CP_4643_elements(69), 
          phi_update_ack => convolve_CP_4643_elements(70), 
          phi_mux_ack => convolve_CP_4643_elements(75), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1926_phi_seq_4942_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4643_elements(92);
      convolve_CP_4643_elements(95)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4643_elements(95);
      convolve_CP_4643_elements(96)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4643_elements(97);
      convolve_CP_4643_elements(93) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4643_elements(90);
      convolve_CP_4643_elements(99)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4643_elements(101);
      convolve_CP_4643_elements(100)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4643_elements(102);
      convolve_CP_4643_elements(91) <= phi_mux_reqs(1);
      phi_stmt_1926_phi_seq_4942 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1926_phi_seq_4942") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4643_elements(86), 
          phi_sample_ack => convolve_CP_4643_elements(87), 
          phi_update_req => convolve_CP_4643_elements(88), 
          phi_update_ack => convolve_CP_4643_elements(89), 
          phi_mux_ack => convolve_CP_4643_elements(94), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1932_phi_seq_4986_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4643_elements(111);
      convolve_CP_4643_elements(114)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4643_elements(114);
      convolve_CP_4643_elements(115)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4643_elements(116);
      convolve_CP_4643_elements(112) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4643_elements(109);
      convolve_CP_4643_elements(118)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4643_elements(120);
      convolve_CP_4643_elements(119)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4643_elements(121);
      convolve_CP_4643_elements(110) <= phi_mux_reqs(1);
      phi_stmt_1932_phi_seq_4986 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1932_phi_seq_4986") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4643_elements(105), 
          phi_sample_ack => convolve_CP_4643_elements(106), 
          phi_update_req => convolve_CP_4643_elements(107), 
          phi_update_ack => convolve_CP_4643_elements(108), 
          phi_mux_ack => convolve_CP_4643_elements(113), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_4762_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convolve_CP_4643_elements(21);
        preds(1)  <= convolve_CP_4643_elements(22);
        entry_tmerge_4762 : transition_merge -- 
          generic map(name => " entry_tmerge_4762")
          port map (preds => preds, symbol_out => convolve_CP_4643_elements(23));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_i16_i16_2136_wire : std_logic_vector(15 downto 0);
    signal ADD_i16_i16_2139_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_2206_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_2226_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_2235_wire : std_logic_vector(15 downto 0);
    signal ADD_u2_u2_2215_wire : std_logic_vector(1 downto 0);
    signal AND_u1_u1_2172_wire : std_logic_vector(0 downto 0);
    signal EQ_u16_u1_1941_wire : std_logic_vector(0 downto 0);
    signal EQ_u16_u1_2043_wire : std_logic_vector(0 downto 0);
    signal EQ_u16_u1_2046_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1944_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2150_wire : std_logic_vector(0 downto 0);
    signal MUL_i16_i16_2115_wire : std_logic_vector(15 downto 0);
    signal MUL_i16_i16_2121_wire : std_logic_vector(15 downto 0);
    signal MUL_i16_i16_2127_wire : std_logic_vector(15 downto 0);
    signal MUX_2216_wire : std_logic_vector(1 downto 0);
    signal MUX_2227_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_2274_wire : std_logic_vector(0 downto 0);
    signal RPIPE_num_out_pipe_1894_wire : std_logic_vector(15 downto 0);
    signal RPIPE_num_out_pipe_1899_wire : std_logic_vector(15 downto 0);
    signal RPIPE_size_pipe_1904_wire : std_logic_vector(15 downto 0);
    signal UGT_u2_u1_2004_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_2001_wire : std_logic_vector(0 downto 0);
    signal acc_1910 : std_logic_vector(15 downto 0);
    signal acc_2059_delayed_1_0_2132 : std_logic_vector(15 downto 0);
    signal acc_val_2141 : std_logic_vector(15 downto 0);
    signal acc_val_dn_2255 : std_logic_vector(7 downto 0);
    signal acc_val_up_2251 : std_logic_vector(7 downto 0);
    signal all_done_flag_2179 : std_logic_vector(0 downto 0);
    signal chl_1932 : std_logic_vector(15 downto 0);
    signal chl_done_2146 : std_logic_vector(0 downto 0);
    signal col_1921 : std_logic_vector(15 downto 0);
    signal col_done_2158 : std_logic_vector(0 downto 0);
    signal iread1_1979 : std_logic_vector(15 downto 0);
    signal iread2_1988 : std_logic_vector(15 downto 0);
    signal iread3_1997 : std_logic_vector(15 downto 0);
    signal ival1_2031 : std_logic_vector(15 downto 0);
    signal ival2_2035 : std_logic_vector(15 downto 0);
    signal ival3_2039 : std_logic_vector(15 downto 0);
    signal konst_1895_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1900_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1905_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1940_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1943_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2003_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2042_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2045_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2149_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2203_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2205_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2212_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2214_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2223_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2225_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2234_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2244_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2276_wire_constant : std_logic_vector(7 downto 0);
    signal kread1_2081 : std_logic_vector(15 downto 0);
    signal kread2_2090 : std_logic_vector(15 downto 0);
    signal kread3_2099 : std_logic_vector(15 downto 0);
    signal kval1_2103 : std_logic_vector(15 downto 0);
    signal kval2_2107 : std_logic_vector(15 downto 0);
    signal kval3_2111 : std_logic_vector(15 downto 0);
    signal mul_val1_2117 : std_logic_vector(15 downto 0);
    signal mul_val2_2123 : std_logic_vector(15 downto 0);
    signal mul_val3_2129 : std_logic_vector(15 downto 0);
    signal n_chl_2208 : std_logic_vector(15 downto 0);
    signal n_chl_2208_1936_buffered : std_logic_vector(15 downto 0);
    signal n_col_2230 : std_logic_vector(15 downto 0);
    signal n_col_2230_1925_buffered : std_logic_vector(15 downto 0);
    signal n_num_2219 : std_logic_vector(1 downto 0);
    signal n_num_2219_1931_buffered : std_logic_vector(1 downto 0);
    signal n_row_2238 : std_logic_vector(15 downto 0);
    signal n_row_2238_1920_buffered : std_logic_vector(15 downto 0);
    signal nacc_2247 : std_logic_vector(15 downto 0);
    signal nacc_2247_1915_buffered : std_logic_vector(15 downto 0);
    signal num_1926 : std_logic_vector(1 downto 0);
    signal num_chl_1907 : std_logic_vector(15 downto 0);
    signal num_col_1902 : std_logic_vector(15 downto 0);
    signal num_done_2153 : std_logic_vector(0 downto 0);
    signal num_done_2156_delayed_1_0_2241 : std_logic_vector(0 downto 0);
    signal num_done_2169_delayed_2_0_2258 : std_logic_vector(0 downto 0);
    signal num_done_2174_delayed_2_0_2266 : std_logic_vector(0 downto 0);
    signal num_row_1897 : std_logic_vector(15 downto 0);
    signal out_done_flag_2168 : std_logic_vector(0 downto 0);
    signal read_ip_1927_delayed_1_0_1973 : std_logic_vector(0 downto 0);
    signal read_ip_1933_delayed_1_0_1982 : std_logic_vector(0 downto 0);
    signal read_ip_1939_delayed_1_0_1991 : std_logic_vector(0 downto 0);
    signal read_ip_1946 : std_logic_vector(0 downto 0);
    signal read_k_2011_delayed_1_0_2075 : std_logic_vector(0 downto 0);
    signal read_k_2017_delayed_1_0_2084 : std_logic_vector(0 downto 0);
    signal read_k_2023_delayed_1_0_2093 : std_logic_vector(0 downto 0);
    signal read_k_2048 : std_logic_vector(0 downto 0);
    signal row_1916 : std_logic_vector(15 downto 0);
    signal row_done_2163 : std_logic_vector(0 downto 0);
    signal store_kernel_2105_delayed_1_0_2182 : std_logic_vector(0 downto 0);
    signal store_kernel_2109_delayed_1_0_2189 : std_logic_vector(0 downto 0);
    signal store_kernel_2113_delayed_1_0_2196 : std_logic_vector(0 downto 0);
    signal store_kernel_2174 : std_logic_vector(0 downto 0);
    signal temp1_1_1962 : std_logic_vector(15 downto 0);
    signal temp1_2_1966 : std_logic_vector(15 downto 0);
    signal temp1_3_1970 : std_logic_vector(15 downto 0);
    signal temp2_1_1950 : std_logic_vector(15 downto 0);
    signal temp2_2_1954 : std_logic_vector(15 downto 0);
    signal temp2_3_1958 : std_logic_vector(15 downto 0);
    signal tempk1_1_2052 : std_logic_vector(15 downto 0);
    signal tempk1_2_2056 : std_logic_vector(15 downto 0);
    signal tempk1_3_2060 : std_logic_vector(15 downto 0);
    signal tempk2_1_2064 : std_logic_vector(15 downto 0);
    signal tempk2_2_2068 : std_logic_vector(15 downto 0);
    signal tempk2_3_2072 : std_logic_vector(15 downto 0);
    signal type_cast_1914_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1919_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1924_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1930_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_1935_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2262_wire : std_logic_vector(7 downto 0);
    signal type_cast_2270_wire : std_logic_vector(7 downto 0);
    signal write_input_1953_delayed_1_0_2009 : std_logic_vector(0 downto 0);
    signal write_input_1957_delayed_1_0_2016 : std_logic_vector(0 downto 0);
    signal write_input_1961_delayed_1_0_2023 : std_logic_vector(0 downto 0);
    signal write_input_2006 : std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip1
    signal xxconvolvexxconv_ip1_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip1_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip1_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip1
    signal xxconvolvexxconv_ip1_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip1_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip1_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip2
    signal xxconvolvexxconv_ip2_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip2_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip2_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip2
    signal xxconvolvexxconv_ip2_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip2_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip2_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip3
    signal xxconvolvexxconv_ip3_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip3_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip3_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip3
    signal xxconvolvexxconv_ip3_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_ip3_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip3_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_k1
    signal xxconvolvexxconv_k1_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k1_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k1_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_k1
    signal xxconvolvexxconv_k1_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k1_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k1_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_k2
    signal xxconvolvexxconv_k2_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k2_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k2_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_k2
    signal xxconvolvexxconv_k2_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k2_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k2_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_k3
    signal xxconvolvexxconv_k3_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k3_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k3_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_k3
    signal xxconvolvexxconv_k3_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxconvolvexxconv_k3_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k3_pipe_read_ack: std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_1895_wire_constant <= "0000000000000001";
    konst_1900_wire_constant <= "0000000000000001";
    konst_1905_wire_constant <= "0000000000000001";
    konst_1940_wire_constant <= "0000000000000000";
    konst_1943_wire_constant <= "10";
    konst_2003_wire_constant <= "00";
    konst_2042_wire_constant <= "0000000000000000";
    konst_2045_wire_constant <= "0000000000000000";
    konst_2149_wire_constant <= "10";
    konst_2203_wire_constant <= "0000000000000000";
    konst_2205_wire_constant <= "0000000000000001";
    konst_2212_wire_constant <= "00";
    konst_2214_wire_constant <= "01";
    konst_2223_wire_constant <= "0000000000000000";
    konst_2225_wire_constant <= "0000000000000001";
    konst_2234_wire_constant <= "0000000000000001";
    konst_2244_wire_constant <= "0000000000000000";
    konst_2276_wire_constant <= "00000001";
    type_cast_1914_wire_constant <= "0000000000000000";
    type_cast_1919_wire_constant <= "0000000000000000";
    type_cast_1924_wire_constant <= "0000000000000000";
    type_cast_1930_wire_constant <= "00";
    type_cast_1935_wire_constant <= "0000000000000000";
    phi_stmt_1910: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1914_wire_constant & nacc_2247_1915_buffered;
      req <= phi_stmt_1910_req_0 & phi_stmt_1910_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1910",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1910_ack_0,
          idata => idata,
          odata => acc_1910,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1910
    phi_stmt_1916: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1919_wire_constant & n_row_2238_1920_buffered;
      req <= phi_stmt_1916_req_0 & phi_stmt_1916_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1916",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1916_ack_0,
          idata => idata,
          odata => row_1916,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1916
    phi_stmt_1921: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1924_wire_constant & n_col_2230_1925_buffered;
      req <= phi_stmt_1921_req_0 & phi_stmt_1921_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1921",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1921_ack_0,
          idata => idata,
          odata => col_1921,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1921
    phi_stmt_1926: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1930_wire_constant & n_num_2219_1931_buffered;
      req <= phi_stmt_1926_req_0 & phi_stmt_1926_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1926",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1926_ack_0,
          idata => idata,
          odata => num_1926,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1926
    phi_stmt_1932: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1935_wire_constant & n_chl_2208_1936_buffered;
      req <= phi_stmt_1932_req_0 & phi_stmt_1932_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1932",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1932_ack_0,
          idata => idata,
          odata => chl_1932,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1932
    -- flow-through select operator MUX_1978_inst
    iread1_1979 <= temp2_1_1950 when (read_ip_1927_delayed_1_0_1973(0) /=  '0') else temp1_1_1962;
    -- flow-through select operator MUX_1987_inst
    iread2_1988 <= temp2_2_1954 when (read_ip_1933_delayed_1_0_1982(0) /=  '0') else temp1_2_1966;
    -- flow-through select operator MUX_1996_inst
    iread3_1997 <= temp2_3_1958 when (read_ip_1939_delayed_1_0_1991(0) /=  '0') else temp1_3_1970;
    -- flow-through select operator MUX_2080_inst
    kread1_2081 <= tempk1_1_2052 when (read_k_2011_delayed_1_0_2075(0) /=  '0') else tempk2_1_2064;
    -- flow-through select operator MUX_2089_inst
    kread2_2090 <= tempk1_2_2056 when (read_k_2017_delayed_1_0_2084(0) /=  '0') else tempk2_2_2068;
    -- flow-through select operator MUX_2098_inst
    kread3_2099 <= tempk1_3_2060 when (read_k_2023_delayed_1_0_2093(0) /=  '0') else tempk2_3_2072;
    -- flow-through select operator MUX_2207_inst
    n_chl_2208 <= konst_2203_wire_constant when (chl_done_2146(0) /=  '0') else ADD_u16_u16_2206_wire;
    -- flow-through select operator MUX_2216_inst
    MUX_2216_wire <= konst_2212_wire_constant when (num_done_2153(0) /=  '0') else ADD_u2_u2_2215_wire;
    -- flow-through select operator MUX_2218_inst
    n_num_2219 <= MUX_2216_wire when (chl_done_2146(0) /=  '0') else num_1926;
    -- flow-through select operator MUX_2227_inst
    MUX_2227_wire <= konst_2223_wire_constant when (col_done_2158(0) /=  '0') else ADD_u16_u16_2226_wire;
    -- flow-through select operator MUX_2229_inst
    n_col_2230 <= MUX_2227_wire when (num_done_2153(0) /=  '0') else col_1921;
    -- flow-through select operator MUX_2237_inst
    n_row_2238 <= ADD_u16_u16_2235_wire when (row_done_2163(0) /=  '0') else row_1916;
    -- flow-through select operator MUX_2246_inst
    nacc_2247 <= konst_2244_wire_constant when (num_done_2156_delayed_1_0_2241(0) /=  '0') else acc_val_2141;
    slice_2250_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2250_inst_req_0;
      slice_2250_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2250_inst_req_1;
      slice_2250_inst_ack_1<= update_ack(0);
      slice_2250_inst: SliceSplitProtocol generic map(name => "slice_2250_inst", in_data_width => 16, high_index => 15, low_index => 8, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => acc_val_2141, dout => acc_val_up_2251, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2254_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2254_inst_req_0;
      slice_2254_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2254_inst_req_1;
      slice_2254_inst_ack_1<= update_ack(0);
      slice_2254_inst: SliceSplitProtocol generic map(name => "slice_2254_inst", in_data_width => 16, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => acc_val_2141, dout => acc_val_dn_2255, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_acc_2059_delayed_1_0_2130_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_acc_2059_delayed_1_0_2130_inst_req_0;
      W_acc_2059_delayed_1_0_2130_inst_ack_0<= wack(0);
      rreq(0) <= W_acc_2059_delayed_1_0_2130_inst_req_1;
      W_acc_2059_delayed_1_0_2130_inst_ack_1<= rack(0);
      W_acc_2059_delayed_1_0_2130_inst : InterlockBuffer generic map ( -- 
        name => "W_acc_2059_delayed_1_0_2130_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_1910,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => acc_2059_delayed_1_0_2132,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_2156_delayed_1_0_2239_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_2156_delayed_1_0_2239_inst_req_0;
      W_num_done_2156_delayed_1_0_2239_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_2156_delayed_1_0_2239_inst_req_1;
      W_num_done_2156_delayed_1_0_2239_inst_ack_1<= rack(0);
      W_num_done_2156_delayed_1_0_2239_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_2156_delayed_1_0_2239_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_2153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_2156_delayed_1_0_2241,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_2169_delayed_2_0_2256_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_2169_delayed_2_0_2256_inst_req_0;
      W_num_done_2169_delayed_2_0_2256_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_2169_delayed_2_0_2256_inst_req_1;
      W_num_done_2169_delayed_2_0_2256_inst_ack_1<= rack(0);
      W_num_done_2169_delayed_2_0_2256_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_2169_delayed_2_0_2256_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_2153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_2169_delayed_2_0_2258,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_2174_delayed_2_0_2264_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_2174_delayed_2_0_2264_inst_req_0;
      W_num_done_2174_delayed_2_0_2264_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_2174_delayed_2_0_2264_inst_req_1;
      W_num_done_2174_delayed_2_0_2264_inst_ack_1<= rack(0);
      W_num_done_2174_delayed_2_0_2264_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_2174_delayed_2_0_2264_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_2153,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_2174_delayed_2_0_2266,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_1927_delayed_1_0_1971_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_1927_delayed_1_0_1971_inst_req_0;
      W_read_ip_1927_delayed_1_0_1971_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_1927_delayed_1_0_1971_inst_req_1;
      W_read_ip_1927_delayed_1_0_1971_inst_ack_1<= rack(0);
      W_read_ip_1927_delayed_1_0_1971_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_1927_delayed_1_0_1971_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_1946,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_1927_delayed_1_0_1973,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_1933_delayed_1_0_1980_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_1933_delayed_1_0_1980_inst_req_0;
      W_read_ip_1933_delayed_1_0_1980_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_1933_delayed_1_0_1980_inst_req_1;
      W_read_ip_1933_delayed_1_0_1980_inst_ack_1<= rack(0);
      W_read_ip_1933_delayed_1_0_1980_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_1933_delayed_1_0_1980_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_1946,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_1933_delayed_1_0_1982,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_1939_delayed_1_0_1989_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_1939_delayed_1_0_1989_inst_req_0;
      W_read_ip_1939_delayed_1_0_1989_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_1939_delayed_1_0_1989_inst_req_1;
      W_read_ip_1939_delayed_1_0_1989_inst_ack_1<= rack(0);
      W_read_ip_1939_delayed_1_0_1989_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_1939_delayed_1_0_1989_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_1946,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_1939_delayed_1_0_1991,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_k_2011_delayed_1_0_2073_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_k_2011_delayed_1_0_2073_inst_req_0;
      W_read_k_2011_delayed_1_0_2073_inst_ack_0<= wack(0);
      rreq(0) <= W_read_k_2011_delayed_1_0_2073_inst_req_1;
      W_read_k_2011_delayed_1_0_2073_inst_ack_1<= rack(0);
      W_read_k_2011_delayed_1_0_2073_inst : InterlockBuffer generic map ( -- 
        name => "W_read_k_2011_delayed_1_0_2073_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_k_2048,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_k_2011_delayed_1_0_2075,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_k_2017_delayed_1_0_2082_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_k_2017_delayed_1_0_2082_inst_req_0;
      W_read_k_2017_delayed_1_0_2082_inst_ack_0<= wack(0);
      rreq(0) <= W_read_k_2017_delayed_1_0_2082_inst_req_1;
      W_read_k_2017_delayed_1_0_2082_inst_ack_1<= rack(0);
      W_read_k_2017_delayed_1_0_2082_inst : InterlockBuffer generic map ( -- 
        name => "W_read_k_2017_delayed_1_0_2082_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_k_2048,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_k_2017_delayed_1_0_2084,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_k_2023_delayed_1_0_2091_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_k_2023_delayed_1_0_2091_inst_req_0;
      W_read_k_2023_delayed_1_0_2091_inst_ack_0<= wack(0);
      rreq(0) <= W_read_k_2023_delayed_1_0_2091_inst_req_1;
      W_read_k_2023_delayed_1_0_2091_inst_ack_1<= rack(0);
      W_read_k_2023_delayed_1_0_2091_inst : InterlockBuffer generic map ( -- 
        name => "W_read_k_2023_delayed_1_0_2091_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_k_2048,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_k_2023_delayed_1_0_2093,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_store_kernel_2105_delayed_1_0_2180_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_store_kernel_2105_delayed_1_0_2180_inst_req_0;
      W_store_kernel_2105_delayed_1_0_2180_inst_ack_0<= wack(0);
      rreq(0) <= W_store_kernel_2105_delayed_1_0_2180_inst_req_1;
      W_store_kernel_2105_delayed_1_0_2180_inst_ack_1<= rack(0);
      W_store_kernel_2105_delayed_1_0_2180_inst : InterlockBuffer generic map ( -- 
        name => "W_store_kernel_2105_delayed_1_0_2180_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => store_kernel_2174,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => store_kernel_2105_delayed_1_0_2182,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_store_kernel_2109_delayed_1_0_2187_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_store_kernel_2109_delayed_1_0_2187_inst_req_0;
      W_store_kernel_2109_delayed_1_0_2187_inst_ack_0<= wack(0);
      rreq(0) <= W_store_kernel_2109_delayed_1_0_2187_inst_req_1;
      W_store_kernel_2109_delayed_1_0_2187_inst_ack_1<= rack(0);
      W_store_kernel_2109_delayed_1_0_2187_inst : InterlockBuffer generic map ( -- 
        name => "W_store_kernel_2109_delayed_1_0_2187_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => store_kernel_2174,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => store_kernel_2109_delayed_1_0_2189,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_store_kernel_2113_delayed_1_0_2194_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_store_kernel_2113_delayed_1_0_2194_inst_req_0;
      W_store_kernel_2113_delayed_1_0_2194_inst_ack_0<= wack(0);
      rreq(0) <= W_store_kernel_2113_delayed_1_0_2194_inst_req_1;
      W_store_kernel_2113_delayed_1_0_2194_inst_ack_1<= rack(0);
      W_store_kernel_2113_delayed_1_0_2194_inst : InterlockBuffer generic map ( -- 
        name => "W_store_kernel_2113_delayed_1_0_2194_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => store_kernel_2174,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => store_kernel_2113_delayed_1_0_2196,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_1953_delayed_1_0_2007_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_1953_delayed_1_0_2007_inst_req_0;
      W_write_input_1953_delayed_1_0_2007_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_1953_delayed_1_0_2007_inst_req_1;
      W_write_input_1953_delayed_1_0_2007_inst_ack_1<= rack(0);
      W_write_input_1953_delayed_1_0_2007_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_1953_delayed_1_0_2007_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_2006,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_1953_delayed_1_0_2009,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_1957_delayed_1_0_2014_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_1957_delayed_1_0_2014_inst_req_0;
      W_write_input_1957_delayed_1_0_2014_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_1957_delayed_1_0_2014_inst_req_1;
      W_write_input_1957_delayed_1_0_2014_inst_ack_1<= rack(0);
      W_write_input_1957_delayed_1_0_2014_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_1957_delayed_1_0_2014_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_2006,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_1957_delayed_1_0_2016,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_1961_delayed_1_0_2021_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_1961_delayed_1_0_2021_inst_req_0;
      W_write_input_1961_delayed_1_0_2021_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_1961_delayed_1_0_2021_inst_req_1;
      W_write_input_1961_delayed_1_0_2021_inst_ack_1<= rack(0);
      W_write_input_1961_delayed_1_0_2021_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_1961_delayed_1_0_2021_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_2006,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_1961_delayed_1_0_2023,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_chl_2208_1936_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_chl_2208_1936_buf_req_0;
      n_chl_2208_1936_buf_ack_0<= wack(0);
      rreq(0) <= n_chl_2208_1936_buf_req_1;
      n_chl_2208_1936_buf_ack_1<= rack(0);
      n_chl_2208_1936_buf : InterlockBuffer generic map ( -- 
        name => "n_chl_2208_1936_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_chl_2208,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_chl_2208_1936_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_col_2230_1925_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_2230_1925_buf_req_0;
      n_col_2230_1925_buf_ack_0<= wack(0);
      rreq(0) <= n_col_2230_1925_buf_req_1;
      n_col_2230_1925_buf_ack_1<= rack(0);
      n_col_2230_1925_buf : InterlockBuffer generic map ( -- 
        name => "n_col_2230_1925_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_2230,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_2230_1925_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_num_2219_1931_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_num_2219_1931_buf_req_0;
      n_num_2219_1931_buf_ack_0<= wack(0);
      rreq(0) <= n_num_2219_1931_buf_req_1;
      n_num_2219_1931_buf_ack_1<= rack(0);
      n_num_2219_1931_buf : InterlockBuffer generic map ( -- 
        name => "n_num_2219_1931_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_num_2219,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_num_2219_1931_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row_2238_1920_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row_2238_1920_buf_req_0;
      n_row_2238_1920_buf_ack_0<= wack(0);
      rreq(0) <= n_row_2238_1920_buf_req_1;
      n_row_2238_1920_buf_ack_1<= rack(0);
      n_row_2238_1920_buf : InterlockBuffer generic map ( -- 
        name => "n_row_2238_1920_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row_2238,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row_2238_1920_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nacc_2247_1915_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nacc_2247_1915_buf_req_0;
      nacc_2247_1915_buf_ack_0<= wack(0);
      rreq(0) <= nacc_2247_1915_buf_req_1;
      nacc_2247_1915_buf_ack_1<= rack(0);
      nacc_2247_1915_buf : InterlockBuffer generic map ( -- 
        name => "nacc_2247_1915_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nacc_2247,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nacc_2247_1915_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2030_inst
    process(iread1_1979) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread1_1979(15 downto 0);
      ival1_2031 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2034_inst
    process(iread2_1988) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread2_1988(15 downto 0);
      ival2_2035 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2038_inst
    process(iread3_1997) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread3_1997(15 downto 0);
      ival3_2039 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2102_inst
    process(kread1_2081) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread1_2081(15 downto 0);
      kval1_2103 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2106_inst
    process(kread2_2090) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread2_2090(15 downto 0);
      kval2_2107 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2110_inst
    process(kread3_2099) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread3_2099(15 downto 0);
      kval3_2111 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2116_inst
    process(MUL_i16_i16_2115_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_i16_i16_2115_wire(15 downto 0);
      mul_val1_2117 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2122_inst
    process(MUL_i16_i16_2121_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_i16_i16_2121_wire(15 downto 0);
      mul_val2_2123 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2128_inst
    process(MUL_i16_i16_2127_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_i16_i16_2127_wire(15 downto 0);
      mul_val3_2129 <= tmp_var; -- 
    end process;
    type_cast_2262_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_2262_inst_req_0;
      type_cast_2262_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_2262_inst_req_1;
      type_cast_2262_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  num_done_2169_delayed_2_0_2258(0);
      type_cast_2262_inst_gI: SplitGuardInterface generic map(name => "type_cast_2262_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_2262_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2262_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val_up_2251,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2262_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2270_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_2270_inst_req_0;
      type_cast_2270_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_2270_inst_req_1;
      type_cast_2270_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  num_done_2174_delayed_2_0_2266(0);
      type_cast_2270_inst_gI: SplitGuardInterface generic map(name => "type_cast_2270_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_2270_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2270_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val_dn_2255,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2270_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1908_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_2274_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1908_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1908_branch_req_0,
          ack0 => do_while_stmt_1908_branch_ack_0,
          ack1 => do_while_stmt_1908_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_i16_i16_2136_inst
    process(acc_2059_delayed_1_0_2132, mul_val1_2117) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(acc_2059_delayed_1_0_2132, mul_val1_2117, tmp_var);
      ADD_i16_i16_2136_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i16_i16_2139_inst
    process(mul_val2_2123, mul_val3_2129) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val2_2123, mul_val3_2129, tmp_var);
      ADD_i16_i16_2139_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i16_i16_2140_inst
    process(ADD_i16_i16_2136_wire, ADD_i16_i16_2139_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i16_i16_2136_wire, ADD_i16_i16_2139_wire, tmp_var);
      acc_val_2141 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2206_inst
    process(chl_1932) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(chl_1932, konst_2205_wire_constant, tmp_var);
      ADD_u16_u16_2206_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2226_inst
    process(col_1921) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_1921, konst_2225_wire_constant, tmp_var);
      ADD_u16_u16_2226_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2235_inst
    process(row_1916) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row_1916, konst_2234_wire_constant, tmp_var);
      ADD_u16_u16_2235_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u2_u2_2215_inst
    process(num_1926) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_1926, konst_2214_wire_constant, tmp_var);
      ADD_u2_u2_2215_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2005_inst
    process(ULT_u16_u1_2001_wire, UGT_u2_u1_2004_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ULT_u16_u1_2001_wire, UGT_u2_u1_2004_wire, tmp_var);
      write_input_2006 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2047_inst
    process(EQ_u16_u1_2043_wire, EQ_u16_u1_2046_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u16_u1_2043_wire, EQ_u16_u1_2046_wire, tmp_var);
      read_k_2048 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2152_inst
    process(EQ_u2_u1_2150_wire, chl_done_2146) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_2150_wire, chl_done_2146, tmp_var);
      num_done_2153 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2162_inst
    process(col_done_2158, num_done_2153) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(col_done_2158, num_done_2153, tmp_var);
      row_done_2163 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2172_inst
    process(out_done_flag_2168, col_done_2158) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_2168, col_done_2158, tmp_var);
      AND_u1_u1_2172_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2178_inst
    process(out_done_flag_2168, row_done_2163) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_2168, row_done_2163, tmp_var);
      all_done_flag_2179 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1941_inst
    process(col_1921) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_1921, konst_1940_wire_constant, tmp_var);
      EQ_u16_u1_1941_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2043_inst
    process(col_1921) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_1921, konst_2042_wire_constant, tmp_var);
      EQ_u16_u1_2043_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2046_inst
    process(row_1916) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(row_1916, konst_2045_wire_constant, tmp_var);
      EQ_u16_u1_2046_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2145_inst
    process(chl_1932, num_chl_1907) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(chl_1932, num_chl_1907, tmp_var);
      chl_done_2146 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2157_inst
    process(col_1921, num_col_1902) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_1921, num_col_1902, tmp_var);
      col_done_2158 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2167_inst
    process(row_1916, num_row_1897) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(row_1916, num_row_1897, tmp_var);
      out_done_flag_2168 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1944_inst
    process(num_1926) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_1926, konst_1943_wire_constant, tmp_var);
      EQ_u2_u1_1944_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_2150_inst
    process(num_1926) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_1926, konst_2149_wire_constant, tmp_var);
      EQ_u2_u1_2150_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_2115_inst
    process(kval1_2103, ival1_2031) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval1_2103, ival1_2031, tmp_var);
      MUL_i16_i16_2115_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_2121_inst
    process(kval2_2107, ival2_2035) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval2_2107, ival2_2035, tmp_var);
      MUL_i16_i16_2121_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_2127_inst
    process(kval3_2111, ival3_2039) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval3_2111, ival3_2039, tmp_var);
      MUL_i16_i16_2127_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_2173_inst
    process(AND_u1_u1_2172_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", AND_u1_u1_2172_wire, tmp_var);
      store_kernel_2174 <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2274_inst
    process(all_done_flag_2179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", all_done_flag_2179, tmp_var);
      NOT_u1_u1_2274_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1945_inst
    process(EQ_u16_u1_1941_wire, EQ_u2_u1_1944_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u16_u1_1941_wire, EQ_u2_u1_1944_wire, tmp_var);
      read_ip_1946 <= tmp_var; --
    end process;
    -- shared split operator group (27) : SUB_u16_u16_1896_inst 
    ApIntSub_group_27: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_num_out_pipe_1894_wire;
      num_row_1897 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_1896_inst_req_0;
      SUB_u16_u16_1896_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_1896_inst_req_1;
      SUB_u16_u16_1896_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_27_gI: SplitGuardInterface generic map(name => "ApIntSub_group_27_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_27",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : SUB_u16_u16_1901_inst 
    ApIntSub_group_28: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_num_out_pipe_1899_wire;
      num_col_1902 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_1901_inst_req_0;
      SUB_u16_u16_1901_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_1901_inst_req_1;
      SUB_u16_u16_1901_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_28_gI: SplitGuardInterface generic map(name => "ApIntSub_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : SUB_u16_u16_1906_inst 
    ApIntSub_group_29: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_size_pipe_1904_wire;
      num_chl_1907 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_1906_inst_req_0;
      SUB_u16_u16_1906_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_1906_inst_req_1;
      SUB_u16_u16_1906_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_29_gI: SplitGuardInterface generic map(name => "ApIntSub_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- binary operator UGT_u2_u1_2004_inst
    process(num_1926) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_1926, konst_2003_wire_constant, tmp_var);
      UGT_u2_u1_2004_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_2001_inst
    process(col_1921, num_col_1902) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(col_1921, num_col_1902, tmp_var);
      ULT_u16_u1_2001_wire <= tmp_var; --
    end process;
    xxconvolvexxconv_ip1_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip1",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip1_pipe_read_req,
        read_ack => xxconvolvexxconv_ip1_pipe_read_ack,
        read_data => xxconvolvexxconv_ip1_pipe_read_data,
        write_req => xxconvolvexxconv_ip1_pipe_write_req,
        write_ack => xxconvolvexxconv_ip1_pipe_write_ack,
        write_data => xxconvolvexxconv_ip1_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_ip2_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip2",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip2_pipe_read_req,
        read_ack => xxconvolvexxconv_ip2_pipe_read_ack,
        read_data => xxconvolvexxconv_ip2_pipe_read_data,
        write_req => xxconvolvexxconv_ip2_pipe_write_req,
        write_ack => xxconvolvexxconv_ip2_pipe_write_ack,
        write_data => xxconvolvexxconv_ip2_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_ip3_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip3",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip3_pipe_read_req,
        read_ack => xxconvolvexxconv_ip3_pipe_read_ack,
        read_data => xxconvolvexxconv_ip3_pipe_read_data,
        write_req => xxconvolvexxconv_ip3_pipe_write_req,
        write_ack => xxconvolvexxconv_ip3_pipe_write_ack,
        write_data => xxconvolvexxconv_ip3_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_k1_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_k1",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_k1_pipe_read_req,
        read_ack => xxconvolvexxconv_k1_pipe_read_ack,
        read_data => xxconvolvexxconv_k1_pipe_read_data,
        write_req => xxconvolvexxconv_k1_pipe_write_req,
        write_ack => xxconvolvexxconv_k1_pipe_write_ack,
        write_data => xxconvolvexxconv_k1_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_k2_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_k2",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_k2_pipe_read_req,
        read_ack => xxconvolvexxconv_k2_pipe_read_ack,
        read_data => xxconvolvexxconv_k2_pipe_read_data,
        write_req => xxconvolvexxconv_k2_pipe_write_req,
        write_ack => xxconvolvexxconv_k2_pipe_write_ack,
        write_data => xxconvolvexxconv_k2_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_k3_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_k3",
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 400 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_k3_pipe_read_req,
        read_ack => xxconvolvexxconv_k3_pipe_read_ack,
        read_data => xxconvolvexxconv_k3_pipe_read_data,
        write_req => xxconvolvexxconv_k3_pipe_write_req,
        write_ack => xxconvolvexxconv_k3_pipe_write_ack,
        write_data => xxconvolvexxconv_k3_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    -- shared inport operator group (0) : RPIPE_input_pipe1_1949_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe1_1949_inst_req_0;
      RPIPE_input_pipe1_1949_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe1_1949_inst_req_1;
      RPIPE_input_pipe1_1949_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_1946(0);
      temp2_1_1950 <= data_out(15 downto 0);
      input_pipe1_read_0_gI: SplitGuardInterface generic map(name => "input_pipe1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe1_read_0: InputPortRevised -- 
        generic map ( name => "input_pipe1_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe1_pipe_read_req(0),
          oack => input_pipe1_pipe_read_ack(0),
          odata => input_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_input_pipe2_1953_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe2_1953_inst_req_0;
      RPIPE_input_pipe2_1953_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe2_1953_inst_req_1;
      RPIPE_input_pipe2_1953_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_1946(0);
      temp2_2_1954 <= data_out(15 downto 0);
      input_pipe2_read_1_gI: SplitGuardInterface generic map(name => "input_pipe2_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe2_read_1: InputPortRevised -- 
        generic map ( name => "input_pipe2_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe2_pipe_read_req(0),
          oack => input_pipe2_pipe_read_ack(0),
          odata => input_pipe2_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_input_pipe3_1957_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe3_1957_inst_req_0;
      RPIPE_input_pipe3_1957_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe3_1957_inst_req_1;
      RPIPE_input_pipe3_1957_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_1946(0);
      temp2_3_1958 <= data_out(15 downto 0);
      input_pipe3_read_2_gI: SplitGuardInterface generic map(name => "input_pipe3_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe3_read_2: InputPortRevised -- 
        generic map ( name => "input_pipe3_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe3_pipe_read_req(0),
          oack => input_pipe3_pipe_read_ack(0),
          odata => input_pipe3_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_kernel_pipe1_2051_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe1_2051_inst_req_0;
      RPIPE_kernel_pipe1_2051_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe1_2051_inst_req_1;
      RPIPE_kernel_pipe1_2051_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_k_2048(0);
      tempk1_1_2052 <= data_out(15 downto 0);
      kernel_pipe1_read_3_gI: SplitGuardInterface generic map(name => "kernel_pipe1_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_read_3: InputPortRevised -- 
        generic map ( name => "kernel_pipe1_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe1_pipe_read_req(0),
          oack => kernel_pipe1_pipe_read_ack(0),
          odata => kernel_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_kernel_pipe2_2055_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe2_2055_inst_req_0;
      RPIPE_kernel_pipe2_2055_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe2_2055_inst_req_1;
      RPIPE_kernel_pipe2_2055_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_k_2048(0);
      tempk1_2_2056 <= data_out(15 downto 0);
      kernel_pipe2_read_4_gI: SplitGuardInterface generic map(name => "kernel_pipe2_read_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe2_read_4: InputPortRevised -- 
        generic map ( name => "kernel_pipe2_read_4", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe2_pipe_read_req(0),
          oack => kernel_pipe2_pipe_read_ack(0),
          odata => kernel_pipe2_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared inport operator group (5) : RPIPE_kernel_pipe3_2059_inst 
    InportGroup_5: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe3_2059_inst_req_0;
      RPIPE_kernel_pipe3_2059_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe3_2059_inst_req_1;
      RPIPE_kernel_pipe3_2059_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_k_2048(0);
      tempk1_3_2060 <= data_out(15 downto 0);
      kernel_pipe3_read_5_gI: SplitGuardInterface generic map(name => "kernel_pipe3_read_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe3_read_5: InputPortRevised -- 
        generic map ( name => "kernel_pipe3_read_5", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe3_pipe_read_req(0),
          oack => kernel_pipe3_pipe_read_ack(0),
          odata => kernel_pipe3_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 5
    -- shared inport operator group (6) : RPIPE_num_out_pipe_1894_inst RPIPE_num_out_pipe_1899_inst 
    InportGroup_6: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_num_out_pipe_1894_inst_req_0;
      reqL_unguarded(0) <= RPIPE_num_out_pipe_1899_inst_req_0;
      RPIPE_num_out_pipe_1894_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_num_out_pipe_1899_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_num_out_pipe_1894_inst_req_1;
      reqR_unguarded(0) <= RPIPE_num_out_pipe_1899_inst_req_1;
      RPIPE_num_out_pipe_1894_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_num_out_pipe_1899_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      RPIPE_num_out_pipe_1894_wire <= data_out(31 downto 16);
      RPIPE_num_out_pipe_1899_wire <= data_out(15 downto 0);
      num_out_pipe_read_6_gI: SplitGuardInterface generic map(name => "num_out_pipe_read_6_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_read_6: InputPortRevised -- 
        generic map ( name => "num_out_pipe_read_6", data_width => 16,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => num_out_pipe_pipe_read_req(0),
          oack => num_out_pipe_pipe_read_ack(0),
          odata => num_out_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 6
    -- shared inport operator group (7) : RPIPE_size_pipe_1904_inst 
    InportGroup_7: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_size_pipe_1904_inst_req_0;
      RPIPE_size_pipe_1904_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_size_pipe_1904_inst_req_1;
      RPIPE_size_pipe_1904_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_size_pipe_1904_wire <= data_out(15 downto 0);
      size_pipe_read_7_gI: SplitGuardInterface generic map(name => "size_pipe_read_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      size_pipe_read_7: InputPortRevised -- 
        generic map ( name => "size_pipe_read_7", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => size_pipe_pipe_read_req(0),
          oack => size_pipe_pipe_read_ack(0),
          odata => size_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 7
    -- shared inport operator group (8) : RPIPE_xxconvolvexxconv_ip1_1961_inst 
    InportGroup_8: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip1_1961_inst_req_0;
      RPIPE_xxconvolvexxconv_ip1_1961_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip1_1961_inst_req_1;
      RPIPE_xxconvolvexxconv_ip1_1961_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_1946(0);
      temp1_1_1962 <= data_out(15 downto 0);
      xxconvolvexxconv_ip1_read_8_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip1_read_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip1_read_8: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip1_read_8", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip1_pipe_read_req(0),
          oack => xxconvolvexxconv_ip1_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 8
    -- shared inport operator group (9) : RPIPE_xxconvolvexxconv_ip2_1965_inst 
    InportGroup_9: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip2_1965_inst_req_0;
      RPIPE_xxconvolvexxconv_ip2_1965_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip2_1965_inst_req_1;
      RPIPE_xxconvolvexxconv_ip2_1965_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_1946(0);
      temp1_2_1966 <= data_out(15 downto 0);
      xxconvolvexxconv_ip2_read_9_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip2_read_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip2_read_9: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip2_read_9", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip2_pipe_read_req(0),
          oack => xxconvolvexxconv_ip2_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip2_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 9
    -- shared inport operator group (10) : RPIPE_xxconvolvexxconv_ip3_1969_inst 
    InportGroup_10: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip3_1969_inst_req_0;
      RPIPE_xxconvolvexxconv_ip3_1969_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip3_1969_inst_req_1;
      RPIPE_xxconvolvexxconv_ip3_1969_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_1946(0);
      temp1_3_1970 <= data_out(15 downto 0);
      xxconvolvexxconv_ip3_read_10_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip3_read_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip3_read_10: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip3_read_10", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip3_pipe_read_req(0),
          oack => xxconvolvexxconv_ip3_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip3_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 10
    -- shared inport operator group (11) : RPIPE_xxconvolvexxconv_k1_2063_inst 
    InportGroup_11: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_k1_2063_inst_req_0;
      RPIPE_xxconvolvexxconv_k1_2063_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_k1_2063_inst_req_1;
      RPIPE_xxconvolvexxconv_k1_2063_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_k_2048(0);
      tempk2_1_2064 <= data_out(15 downto 0);
      xxconvolvexxconv_k1_read_11_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k1_read_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k1_read_11: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k1_read_11", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_k1_pipe_read_req(0),
          oack => xxconvolvexxconv_k1_pipe_read_ack(0),
          odata => xxconvolvexxconv_k1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 11
    -- shared inport operator group (12) : RPIPE_xxconvolvexxconv_k2_2067_inst 
    InportGroup_12: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_k2_2067_inst_req_0;
      RPIPE_xxconvolvexxconv_k2_2067_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_k2_2067_inst_req_1;
      RPIPE_xxconvolvexxconv_k2_2067_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_k_2048(0);
      tempk2_2_2068 <= data_out(15 downto 0);
      xxconvolvexxconv_k2_read_12_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k2_read_12_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k2_read_12: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k2_read_12", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_k2_pipe_read_req(0),
          oack => xxconvolvexxconv_k2_pipe_read_ack(0),
          odata => xxconvolvexxconv_k2_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 12
    -- shared inport operator group (13) : RPIPE_xxconvolvexxconv_k3_2071_inst 
    InportGroup_13: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_k3_2071_inst_req_0;
      RPIPE_xxconvolvexxconv_k3_2071_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_k3_2071_inst_req_1;
      RPIPE_xxconvolvexxconv_k3_2071_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_k_2048(0);
      tempk2_3_2072 <= data_out(15 downto 0);
      xxconvolvexxconv_k3_read_13_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k3_read_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k3_read_13: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k3_read_13", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_k3_pipe_read_req(0),
          oack => xxconvolvexxconv_k3_pipe_read_ack(0),
          odata => xxconvolvexxconv_k3_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 13
    -- shared outport operator group (0) : WPIPE_input_done_pipe_2275_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_2275_inst_req_0;
      WPIPE_input_done_pipe_2275_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_2275_inst_req_1;
      WPIPE_input_done_pipe_2275_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_2276_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_maxpool_output_pipe_2260_inst WPIPE_maxpool_output_pipe_2268_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_2260_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_2268_inst_req_0;
      WPIPE_maxpool_output_pipe_2260_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_2268_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_2260_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_2268_inst_req_1;
      WPIPE_maxpool_output_pipe_2260_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_2268_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= num_done_2174_delayed_2_0_2266(0);
      guard_vector(1)  <= num_done_2169_delayed_2_0_2258(0);
      data_in <= type_cast_2262_wire & type_cast_2270_wire;
      maxpool_output_pipe_write_1_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 2, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_xxconvolvexxconv_ip1_2011_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip1_2011_inst_req_0;
      WPIPE_xxconvolvexxconv_ip1_2011_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip1_2011_inst_req_1;
      WPIPE_xxconvolvexxconv_ip1_2011_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_1953_delayed_1_0_2009(0);
      data_in <= iread1_1979;
      xxconvolvexxconv_ip1_write_2_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip1_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip1_write_2: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip1_pipe_write_req(0),
          oack => xxconvolvexxconv_ip1_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_xxconvolvexxconv_ip2_2018_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip2_2018_inst_req_0;
      WPIPE_xxconvolvexxconv_ip2_2018_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip2_2018_inst_req_1;
      WPIPE_xxconvolvexxconv_ip2_2018_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_1957_delayed_1_0_2016(0);
      data_in <= iread2_1988;
      xxconvolvexxconv_ip2_write_3_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip2_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip2_write_3: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip2_pipe_write_req(0),
          oack => xxconvolvexxconv_ip2_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_xxconvolvexxconv_ip3_2025_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip3_2025_inst_req_0;
      WPIPE_xxconvolvexxconv_ip3_2025_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip3_2025_inst_req_1;
      WPIPE_xxconvolvexxconv_ip3_2025_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_1961_delayed_1_0_2023(0);
      data_in <= iread3_1997;
      xxconvolvexxconv_ip3_write_4_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip3_write_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip3_write_4: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip3", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip3_pipe_write_req(0),
          oack => xxconvolvexxconv_ip3_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip3_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared outport operator group (5) : WPIPE_xxconvolvexxconv_k1_2184_inst 
    OutportGroup_5: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k1_2184_inst_req_0;
      WPIPE_xxconvolvexxconv_k1_2184_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k1_2184_inst_req_1;
      WPIPE_xxconvolvexxconv_k1_2184_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= store_kernel_2105_delayed_1_0_2182(0);
      data_in <= kread1_2081;
      xxconvolvexxconv_k1_write_5_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k1_write_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k1_write_5: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_k1_pipe_write_req(0),
          oack => xxconvolvexxconv_k1_pipe_write_ack(0),
          odata => xxconvolvexxconv_k1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- shared outport operator group (6) : WPIPE_xxconvolvexxconv_k2_2191_inst 
    OutportGroup_6: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k2_2191_inst_req_0;
      WPIPE_xxconvolvexxconv_k2_2191_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k2_2191_inst_req_1;
      WPIPE_xxconvolvexxconv_k2_2191_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= store_kernel_2109_delayed_1_0_2189(0);
      data_in <= kread2_2090;
      xxconvolvexxconv_k2_write_6_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k2_write_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k2_write_6: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_k2_pipe_write_req(0),
          oack => xxconvolvexxconv_k2_pipe_write_ack(0),
          odata => xxconvolvexxconv_k2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 6
    -- shared outport operator group (7) : WPIPE_xxconvolvexxconv_k3_2198_inst 
    OutportGroup_7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k3_2198_inst_req_0;
      WPIPE_xxconvolvexxconv_k3_2198_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k3_2198_inst_req_1;
      WPIPE_xxconvolvexxconv_k3_2198_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= store_kernel_2113_delayed_1_0_2196(0);
      data_in <= kread3_2099;
      xxconvolvexxconv_k3_write_7_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k3_write_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k3_write_7: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k3", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_k3_pipe_write_req(0),
          oack => xxconvolvexxconv_k3_pipe_write_ack(0),
          odata => xxconvolvexxconv_k3_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 7
    -- 
  end Block; -- data_path
  -- 
end convolve_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity loadKernelChannel is -- 
  generic (tag_length : integer); 
  port ( -- 
    start_add : in  std_logic_vector(63 downto 0);
    num_chl : in  std_logic_vector(15 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
    kernel_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadKernelChannel;
architecture loadKernelChannel_arch of loadKernelChannel is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 80)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal start_add_buffer :  std_logic_vector(63 downto 0);
  signal start_add_update_enable: Boolean;
  signal num_chl_buffer :  std_logic_vector(15 downto 0);
  signal num_chl_update_enable: Boolean;
  -- output port buffer signals
  signal loadKernelChannel_CP_1309_start: Boolean;
  signal loadKernelChannel_CP_1309_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal phi_stmt_447_req_1 : boolean;
  signal ptr_deref_413_load_0_req_0 : boolean;
  signal start_add_449_buf_ack_0 : boolean;
  signal array_obj_ref_408_index_offset_req_0 : boolean;
  signal start_add_449_buf_req_1 : boolean;
  signal ptr_deref_413_load_0_ack_1 : boolean;
  signal ptr_deref_413_load_0_ack_0 : boolean;
  signal nfetch_val_541_453_buf_req_0 : boolean;
  signal phi_stmt_447_ack_0 : boolean;
  signal addr_of_409_final_reg_req_1 : boolean;
  signal phi_stmt_447_req_0 : boolean;
  signal my_fetch_414_454_buf_req_1 : boolean;
  signal do_while_stmt_445_branch_req_0 : boolean;
  signal start_add_449_buf_ack_1 : boolean;
  signal my_fetch_414_454_buf_req_0 : boolean;
  signal RPIPE_input_done_pipe_442_inst_req_1 : boolean;
  signal ptr_deref_413_load_0_req_1 : boolean;
  signal start_add_449_buf_req_0 : boolean;
  signal RPIPE_input_done_pipe_442_inst_ack_0 : boolean;
  signal nmycount_469_450_buf_ack_1 : boolean;
  signal nfetch_val_541_453_buf_ack_1 : boolean;
  signal nfetch_val_541_453_buf_req_1 : boolean;
  signal RPIPE_input_done_pipe_442_inst_req_0 : boolean;
  signal addr_of_409_final_reg_ack_1 : boolean;
  signal phi_stmt_451_req_1 : boolean;
  signal my_fetch_414_454_buf_ack_1 : boolean;
  signal phi_stmt_451_req_0 : boolean;
  signal WPIPE_kernel_pipe1_495_inst_req_0 : boolean;
  signal nmycount_469_450_buf_req_1 : boolean;
  signal nfetch_val_541_453_buf_ack_0 : boolean;
  signal nmycount_469_450_buf_req_0 : boolean;
  signal WPIPE_kernel_pipe3_503_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe3_503_inst_ack_1 : boolean;
  signal phi_stmt_451_ack_0 : boolean;
  signal addr_of_409_final_reg_req_0 : boolean;
  signal WPIPE_kernel_pipe1_495_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe2_499_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe1_495_inst_ack_0 : boolean;
  signal array_obj_ref_408_index_offset_ack_1 : boolean;
  signal nmycount_469_450_buf_ack_0 : boolean;
  signal WPIPE_kernel_pipe2_499_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe3_503_inst_ack_0 : boolean;
  signal my_fetch_414_454_buf_ack_0 : boolean;
  signal WPIPE_kernel_pipe2_499_inst_ack_0 : boolean;
  signal array_obj_ref_408_index_offset_req_1 : boolean;
  signal WPIPE_kernel_pipe1_495_inst_req_1 : boolean;
  signal addr_of_409_final_reg_ack_0 : boolean;
  signal WPIPE_kernel_pipe3_503_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe2_499_inst_ack_1 : boolean;
  signal RPIPE_input_done_pipe_442_inst_ack_1 : boolean;
  signal array_obj_ref_408_index_offset_ack_0 : boolean;
  signal array_obj_ref_519_index_offset_req_0 : boolean;
  signal array_obj_ref_519_index_offset_ack_0 : boolean;
  signal array_obj_ref_519_index_offset_req_1 : boolean;
  signal array_obj_ref_519_index_offset_ack_1 : boolean;
  signal addr_of_520_final_reg_req_0 : boolean;
  signal addr_of_520_final_reg_ack_0 : boolean;
  signal addr_of_520_final_reg_req_1 : boolean;
  signal addr_of_520_final_reg_ack_1 : boolean;
  signal W_fn_486_delayed_7_0_522_inst_req_0 : boolean;
  signal W_fn_486_delayed_7_0_522_inst_ack_0 : boolean;
  signal W_fn_486_delayed_7_0_522_inst_req_1 : boolean;
  signal W_fn_486_delayed_7_0_522_inst_ack_1 : boolean;
  signal ptr_deref_528_load_0_req_0 : boolean;
  signal ptr_deref_528_load_0_ack_0 : boolean;
  signal ptr_deref_528_load_0_req_1 : boolean;
  signal ptr_deref_528_load_0_ack_1 : boolean;
  signal W_fn_492_delayed_13_0_530_inst_req_0 : boolean;
  signal W_fn_492_delayed_13_0_530_inst_ack_0 : boolean;
  signal W_fn_492_delayed_13_0_530_inst_req_1 : boolean;
  signal W_fn_492_delayed_13_0_530_inst_ack_1 : boolean;
  signal W_fetch_val_494_delayed_13_0_533_inst_req_0 : boolean;
  signal W_fetch_val_494_delayed_13_0_533_inst_ack_0 : boolean;
  signal W_fetch_val_494_delayed_13_0_533_inst_req_1 : boolean;
  signal W_fetch_val_494_delayed_13_0_533_inst_ack_1 : boolean;
  signal do_while_stmt_445_branch_ack_0 : boolean;
  signal do_while_stmt_445_branch_ack_1 : boolean;
  signal WPIPE_size_pipe_549_inst_req_0 : boolean;
  signal WPIPE_size_pipe_549_inst_ack_0 : boolean;
  signal WPIPE_size_pipe_549_inst_req_1 : boolean;
  signal WPIPE_size_pipe_549_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadKernelChannel_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 80) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= start_add;
  start_add_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(79 downto 64) <= num_chl;
  num_chl_buffer <= in_buffer_data_out(79 downto 64);
  in_buffer_data_in(tag_length + 79 downto 80) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 79 downto 80);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadKernelChannel_CP_1309_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadKernelChannel_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_1309_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadKernelChannel_CP_1309_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_1309_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadKernelChannel_CP_1309: Block -- control-path 
    signal loadKernelChannel_CP_1309_elements: BooleanArray(98 downto 0);
    -- 
  begin -- 
    loadKernelChannel_CP_1309_elements(0) <= loadKernelChannel_CP_1309_start;
    loadKernelChannel_CP_1309_symbol <= loadKernelChannel_CP_1309_elements(98);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	7 
    -- CP-element group 0:  members (29) 
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/addr_of_409_complete/$entry
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/RPIPE_input_done_pipe_442_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_index_resized_1
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_update_start_
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/RPIPE_input_done_pipe_442_sample_start_
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/addr_of_409_complete/req
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_index_computed_1
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/addr_of_409_update_start_
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Update/$entry
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/RPIPE_input_done_pipe_442_Sample/rr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/$entry
      -- CP-element group 0: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_final_index_sum_regn_Update/$entry
      -- 
    req_1359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(0), ack => addr_of_409_final_reg_req_1); -- 
    req_1339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(0), ack => array_obj_ref_408_index_offset_req_0); -- 
    req_1344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(0), ack => array_obj_ref_408_index_offset_req_1); -- 
    cr_1404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(0), ack => ptr_deref_413_load_0_req_1); -- 
    rr_1418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(0), ack => RPIPE_input_done_pipe_442_inst_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_final_index_sum_regn_sample_complete
      -- CP-element group 1: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_final_index_sum_regn_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_final_index_sum_regn_Sample/ack
      -- 
    ack_1340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_408_index_offset_ack_0, ack => loadKernelChannel_CP_1309_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_offset_calculated
      -- CP-element group 2: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_base_plus_offset/$entry
      -- CP-element group 2: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 assign_stmt_398_to_assign_stmt_443/addr_of_409_request/$entry
      -- CP-element group 2: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 assign_stmt_398_to_assign_stmt_443/addr_of_409_sample_start_
      -- CP-element group 2: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_root_address_calculated
      -- CP-element group 2: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_base_plus_offset/$exit
      -- CP-element group 2: 	 assign_stmt_398_to_assign_stmt_443/addr_of_409_request/req
      -- CP-element group 2: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_final_index_sum_regn_Update/ack
      -- CP-element group 2: 	 assign_stmt_398_to_assign_stmt_443/array_obj_ref_408_final_index_sum_regn_Update/$exit
      -- 
    ack_1345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_408_index_offset_ack_1, ack => loadKernelChannel_CP_1309_elements(2)); -- 
    req_1354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(2), ack => addr_of_409_final_reg_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_398_to_assign_stmt_443/addr_of_409_request/$exit
      -- CP-element group 3: 	 assign_stmt_398_to_assign_stmt_443/addr_of_409_sample_completed_
      -- CP-element group 3: 	 assign_stmt_398_to_assign_stmt_443/addr_of_409_request/ack
      -- 
    ack_1355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_409_final_reg_ack_0, ack => loadKernelChannel_CP_1309_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (24) 
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_word_address_calculated
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_base_plus_offset/$entry
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_word_addrgen/root_register_req
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_base_plus_offset/sum_rename_ack
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/addr_of_409_update_completed_
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Sample/word_access_start/word_0/rr
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/addr_of_409_complete/$exit
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_base_plus_offset/$exit
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_base_addr_resize/base_resize_ack
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_base_plus_offset/sum_rename_req
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_sample_start_
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_base_address_calculated
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_root_address_calculated
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/addr_of_409_complete/ack
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Sample/word_access_start/word_0/$entry
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_base_address_resized
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_base_addr_resize/$entry
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_word_addrgen/$entry
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_base_addr_resize/$exit
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_word_addrgen/root_register_ack
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Sample/word_access_start/$entry
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_word_addrgen/$exit
      -- CP-element group 4: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_base_addr_resize/base_resize_req
      -- 
    ack_1360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_409_final_reg_ack_1, ack => loadKernelChannel_CP_1309_elements(4)); -- 
    rr_1393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(4), ack => ptr_deref_413_load_0_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Sample/word_access_start/word_0/ra
      -- CP-element group 5: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Sample/word_access_start/$exit
      -- CP-element group 5: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_sample_completed_
      -- CP-element group 5: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Sample/$exit
      -- 
    ra_1394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_413_load_0_ack_0, ack => loadKernelChannel_CP_1309_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_update_completed_
      -- CP-element group 6: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Update/ptr_deref_413_Merge/merge_ack
      -- CP-element group 6: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Update/ptr_deref_413_Merge/merge_req
      -- CP-element group 6: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Update/ptr_deref_413_Merge/$exit
      -- CP-element group 6: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Update/ptr_deref_413_Merge/$entry
      -- CP-element group 6: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Update/word_access_complete/$exit
      -- CP-element group 6: 	 assign_stmt_398_to_assign_stmt_443/ptr_deref_413_Update/$exit
      -- 
    ca_1405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_413_load_0_ack_1, ack => loadKernelChannel_CP_1309_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_398_to_assign_stmt_443/RPIPE_input_done_pipe_442_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_398_to_assign_stmt_443/RPIPE_input_done_pipe_442_update_start_
      -- CP-element group 7: 	 assign_stmt_398_to_assign_stmt_443/RPIPE_input_done_pipe_442_sample_completed_
      -- CP-element group 7: 	 assign_stmt_398_to_assign_stmt_443/RPIPE_input_done_pipe_442_Update/cr
      -- CP-element group 7: 	 assign_stmt_398_to_assign_stmt_443/RPIPE_input_done_pipe_442_Update/$entry
      -- CP-element group 7: 	 assign_stmt_398_to_assign_stmt_443/RPIPE_input_done_pipe_442_Sample/ra
      -- 
    ra_1419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_442_inst_ack_0, ack => loadKernelChannel_CP_1309_elements(7)); -- 
    cr_1423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(7), ack => RPIPE_input_done_pipe_442_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_398_to_assign_stmt_443/RPIPE_input_done_pipe_442_update_completed_
      -- CP-element group 8: 	 assign_stmt_398_to_assign_stmt_443/RPIPE_input_done_pipe_442_Update/$exit
      -- CP-element group 8: 	 assign_stmt_398_to_assign_stmt_443/RPIPE_input_done_pipe_442_Update/ca
      -- 
    ca_1424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_442_inst_ack_1, ack => loadKernelChannel_CP_1309_elements(8)); -- 
    -- CP-element group 9:  join  transition  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: 	6 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 assign_stmt_398_to_assign_stmt_443/$exit
      -- CP-element group 9: 	 branch_block_stmt_444/do_while_stmt_445__entry__
      -- CP-element group 9: 	 branch_block_stmt_444/branch_block_stmt_444__entry__
      -- CP-element group 9: 	 branch_block_stmt_444/$entry
      -- 
    loadKernelChannel_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 36) := "loadKernelChannel_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(1) & loadKernelChannel_CP_1309_elements(6) & loadKernelChannel_CP_1309_elements(8);
      gj_loadKernelChannel_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  transition  place  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	96 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	97 
    -- CP-element group 10:  members (7) 
      -- CP-element group 10: 	 branch_block_stmt_444/do_while_stmt_445__exit__
      -- CP-element group 10: 	 branch_block_stmt_444/branch_block_stmt_444__exit__
      -- CP-element group 10: 	 branch_block_stmt_444/$exit
      -- CP-element group 10: 	 assign_stmt_551/$entry
      -- CP-element group 10: 	 assign_stmt_551/WPIPE_size_pipe_549_sample_start_
      -- CP-element group 10: 	 assign_stmt_551/WPIPE_size_pipe_549_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_551/WPIPE_size_pipe_549_Sample/req
      -- 
    req_1760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(10), ack => WPIPE_size_pipe_549_inst_req_0); -- 
    loadKernelChannel_CP_1309_elements(10) <= loadKernelChannel_CP_1309_elements(96);
    -- CP-element group 11:  transition  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445__entry__
      -- CP-element group 11: 	 branch_block_stmt_444/do_while_stmt_445/$entry
      -- 
    loadKernelChannel_CP_1309_elements(11) <= loadKernelChannel_CP_1309_elements(9);
    -- CP-element group 12:  merge  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	96 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445__exit__
      -- 
    -- Element group loadKernelChannel_CP_1309_elements(12) is bound as output of CP function.
    -- CP-element group 13:  merge  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	16 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_444/do_while_stmt_445/loop_back
      -- 
    -- Element group loadKernelChannel_CP_1309_elements(13) is bound as output of CP function.
    -- CP-element group 14:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	95 
    -- CP-element group 14: 	94 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_444/do_while_stmt_445/condition_done
      -- CP-element group 14: 	 branch_block_stmt_444/do_while_stmt_445/loop_exit/$entry
      -- CP-element group 14: 	 branch_block_stmt_444/do_while_stmt_445/loop_taken/$entry
      -- 
    loadKernelChannel_CP_1309_elements(14) <= loadKernelChannel_CP_1309_elements(19);
    -- CP-element group 15:  branch  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	93 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_444/do_while_stmt_445/loop_body_done
      -- 
    loadKernelChannel_CP_1309_elements(15) <= loadKernelChannel_CP_1309_elements(93);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	13 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	28 
    -- CP-element group 16: 	47 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/back_edge_to_loop_body
      -- 
    loadKernelChannel_CP_1309_elements(16) <= loadKernelChannel_CP_1309_elements(13);
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	30 
    -- CP-element group 17: 	49 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/first_time_through_loop_body
      -- 
    loadKernelChannel_CP_1309_elements(17) <= loadKernelChannel_CP_1309_elements(11);
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	92 
    -- CP-element group 18: 	24 
    -- CP-element group 18: 	25 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	42 
    -- CP-element group 18: 	70 
    -- CP-element group 18: 	71 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/$entry
      -- CP-element group 18: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/loop_body_start
      -- 
    -- Element group loadKernelChannel_CP_1309_elements(18) is bound as output of CP function.
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	92 
    -- CP-element group 19: 	23 
    -- CP-element group 19: 	27 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/condition_evaluated
      -- 
    condition_evaluated_1446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(19), ack => do_while_stmt_445_branch_req_0); -- 
    loadKernelChannel_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(92) & loadKernelChannel_CP_1309_elements(23) & loadKernelChannel_CP_1309_elements(27);
      gj_loadKernelChannel_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	24 
    -- CP-element group 20: 	41 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	23 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	43 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/aggregated_phi_sample_req
      -- CP-element group 20: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_447_sample_start__ps
      -- 
    loadKernelChannel_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(24) & loadKernelChannel_CP_1309_elements(41) & loadKernelChannel_CP_1309_elements(23);
      gj_loadKernelChannel_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	26 
    -- CP-element group 21: 	44 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	93 
    -- CP-element group 21: 	81 
    -- CP-element group 21: 	85 
    -- CP-element group 21: 	89 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	24 
    -- CP-element group 21: 	41 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_451_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/aggregated_phi_sample_ack
      -- CP-element group 21: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_447_sample_completed_
      -- 
    loadKernelChannel_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(26) & loadKernelChannel_CP_1309_elements(44);
      gj_loadKernelChannel_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	25 
    -- CP-element group 22: 	42 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	45 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/aggregated_phi_update_req
      -- CP-element group 22: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_447_update_start__ps
      -- 
    loadKernelChannel_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(25) & loadKernelChannel_CP_1309_elements(42);
      gj_loadKernelChannel_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	27 
    -- CP-element group 23: 	46 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/aggregated_phi_update_ack
      -- 
    loadKernelChannel_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(27) & loadKernelChannel_CP_1309_elements(46);
      gj_loadKernelChannel_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	20 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_447_sample_start_
      -- 
    loadKernelChannel_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(18) & loadKernelChannel_CP_1309_elements(21);
      gj_loadKernelChannel_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	18 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	27 
    -- CP-element group 25: 	61 
    -- CP-element group 25: 	64 
    -- CP-element group 25: 	67 
    -- CP-element group 25: 	72 
    -- CP-element group 25: 	78 
    -- CP-element group 25: 	86 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	22 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_447_update_start_
      -- 
    loadKernelChannel_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1,6 => 0,7 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(18) & loadKernelChannel_CP_1309_elements(27) & loadKernelChannel_CP_1309_elements(61) & loadKernelChannel_CP_1309_elements(64) & loadKernelChannel_CP_1309_elements(67) & loadKernelChannel_CP_1309_elements(72) & loadKernelChannel_CP_1309_elements(78) & loadKernelChannel_CP_1309_elements(86);
      gj_loadKernelChannel_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	21 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_447_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_1309_elements(26) is bound as output of CP function.
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	19 
    -- CP-element group 27: 	23 
    -- CP-element group 27: 	60 
    -- CP-element group 27: 	63 
    -- CP-element group 27: 	66 
    -- CP-element group 27: 	72 
    -- CP-element group 27: 	76 
    -- CP-element group 27: 	84 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	25 
    -- CP-element group 27:  members (15) 
      -- CP-element group 27: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_447_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_index_resize_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_index_scale_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_index_scale_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_index_resize_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_index_resize_1/index_resize_req
      -- CP-element group 27: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_index_resized_1
      -- CP-element group 27: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_index_resize_1/index_resize_ack
      -- CP-element group 27: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_index_scale_1/scale_rename_req
      -- CP-element group 27: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_index_computed_1
      -- CP-element group 27: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_index_scale_1/scale_rename_ack
      -- CP-element group 27: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_final_index_sum_regn_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_index_scaled_1
      -- CP-element group 27: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_447_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_final_index_sum_regn_Sample/req
      -- 
    req_1626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(27), ack => array_obj_ref_519_index_offset_req_0); -- 
    -- Element group loadKernelChannel_CP_1309_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	16 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_447_loopback_trigger
      -- 
    loadKernelChannel_CP_1309_elements(28) <= loadKernelChannel_CP_1309_elements(16);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_447_loopback_sample_req
      -- CP-element group 29: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_447_loopback_sample_req_ps
      -- 
    phi_stmt_447_loopback_sample_req_1461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_447_loopback_sample_req_1461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(29), ack => phi_stmt_447_req_1); -- 
    -- Element group loadKernelChannel_CP_1309_elements(29) is bound as output of CP function.
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	17 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_447_entry_trigger
      -- 
    loadKernelChannel_CP_1309_elements(30) <= loadKernelChannel_CP_1309_elements(17);
    -- CP-element group 31:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_447_entry_sample_req_ps
      -- CP-element group 31: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_447_entry_sample_req
      -- 
    phi_stmt_447_entry_sample_req_1464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_447_entry_sample_req_1464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(31), ack => phi_stmt_447_req_0); -- 
    -- Element group loadKernelChannel_CP_1309_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_447_phi_mux_ack_ps
      -- CP-element group 32: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_447_phi_mux_ack
      -- 
    phi_stmt_447_phi_mux_ack_1467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_447_ack_0, ack => loadKernelChannel_CP_1309_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_start_add_449_sample_start__ps
      -- CP-element group 33: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_start_add_449_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_start_add_449_Sample/req
      -- CP-element group 33: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_start_add_449_Sample/$entry
      -- 
    req_1480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(33), ack => start_add_449_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1309_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_start_add_449_Update/req
      -- CP-element group 34: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_start_add_449_update_start__ps
      -- CP-element group 34: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_start_add_449_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_start_add_449_update_start_
      -- 
    req_1485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(34), ack => start_add_449_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1309_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_start_add_449_sample_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_start_add_449_Sample/ack
      -- CP-element group 35: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_start_add_449_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_start_add_449_sample_completed_
      -- 
    ack_1481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_449_buf_ack_0, ack => loadKernelChannel_CP_1309_elements(35)); -- 
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_start_add_449_update_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_start_add_449_Update/ack
      -- CP-element group 36: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_start_add_449_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_start_add_449_update_completed_
      -- 
    ack_1486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_449_buf_ack_1, ack => loadKernelChannel_CP_1309_elements(36)); -- 
    -- CP-element group 37:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nmycount_450_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nmycount_450_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nmycount_450_sample_start__ps
      -- CP-element group 37: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nmycount_450_Sample/req
      -- 
    req_1498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(37), ack => nmycount_469_450_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1309_elements(37) is bound as output of CP function.
    -- CP-element group 38:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nmycount_450_update_start_
      -- CP-element group 38: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nmycount_450_update_start__ps
      -- CP-element group 38: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nmycount_450_Update/req
      -- CP-element group 38: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nmycount_450_Update/$entry
      -- 
    req_1503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(38), ack => nmycount_469_450_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1309_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nmycount_450_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nmycount_450_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nmycount_450_sample_completed__ps
      -- CP-element group 39: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nmycount_450_Sample/ack
      -- 
    ack_1499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_469_450_buf_ack_0, ack => loadKernelChannel_CP_1309_elements(39)); -- 
    -- CP-element group 40:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nmycount_450_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nmycount_450_update_completed__ps
      -- CP-element group 40: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nmycount_450_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nmycount_450_Update/ack
      -- 
    ack_1504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_469_450_buf_ack_1, ack => loadKernelChannel_CP_1309_elements(40)); -- 
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	91 
    -- CP-element group 41: 	21 
    -- CP-element group 41: 	83 
    -- CP-element group 41: 	87 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	20 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_451_sample_start_
      -- 
    loadKernelChannel_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(18) & loadKernelChannel_CP_1309_elements(91) & loadKernelChannel_CP_1309_elements(21) & loadKernelChannel_CP_1309_elements(83) & loadKernelChannel_CP_1309_elements(87);
      gj_loadKernelChannel_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	18 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	90 
    -- CP-element group 42: 	46 
    -- CP-element group 42: 	61 
    -- CP-element group 42: 	64 
    -- CP-element group 42: 	67 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	22 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_451_update_start_
      -- 
    loadKernelChannel_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(18) & loadKernelChannel_CP_1309_elements(90) & loadKernelChannel_CP_1309_elements(46) & loadKernelChannel_CP_1309_elements(61) & loadKernelChannel_CP_1309_elements(64) & loadKernelChannel_CP_1309_elements(67);
      gj_loadKernelChannel_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	20 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_451_sample_start__ps
      -- 
    loadKernelChannel_CP_1309_elements(43) <= loadKernelChannel_CP_1309_elements(20);
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	21 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_451_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_1309_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	22 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_451_update_start__ps
      -- 
    loadKernelChannel_CP_1309_elements(45) <= loadKernelChannel_CP_1309_elements(22);
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	23 
    -- CP-element group 46: 	60 
    -- CP-element group 46: 	63 
    -- CP-element group 46: 	66 
    -- CP-element group 46: 	88 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	42 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_451_update_completed__ps
      -- CP-element group 46: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_451_update_completed_
      -- 
    -- Element group loadKernelChannel_CP_1309_elements(46) is bound as output of CP function.
    -- CP-element group 47:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	16 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_451_loopback_trigger
      -- 
    loadKernelChannel_CP_1309_elements(47) <= loadKernelChannel_CP_1309_elements(16);
    -- CP-element group 48:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_451_loopback_sample_req_ps
      -- CP-element group 48: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_451_loopback_sample_req
      -- 
    phi_stmt_451_loopback_sample_req_1515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_451_loopback_sample_req_1515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(48), ack => phi_stmt_451_req_0); -- 
    -- Element group loadKernelChannel_CP_1309_elements(48) is bound as output of CP function.
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	17 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_451_entry_trigger
      -- 
    loadKernelChannel_CP_1309_elements(49) <= loadKernelChannel_CP_1309_elements(17);
    -- CP-element group 50:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_451_entry_sample_req
      -- CP-element group 50: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_451_entry_sample_req_ps
      -- 
    phi_stmt_451_entry_sample_req_1518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_451_entry_sample_req_1518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(50), ack => phi_stmt_451_req_1); -- 
    -- Element group loadKernelChannel_CP_1309_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_451_phi_mux_ack
      -- CP-element group 51: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/phi_stmt_451_phi_mux_ack_ps
      -- 
    phi_stmt_451_phi_mux_ack_1521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_451_ack_0, ack => loadKernelChannel_CP_1309_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nfetch_val_453_Sample/req
      -- CP-element group 52: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nfetch_val_453_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nfetch_val_453_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nfetch_val_453_sample_start__ps
      -- 
    req_1534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(52), ack => nfetch_val_541_453_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1309_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nfetch_val_453_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nfetch_val_453_update_start_
      -- CP-element group 53: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nfetch_val_453_Update/req
      -- CP-element group 53: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nfetch_val_453_Update/$entry
      -- 
    req_1539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(53), ack => nfetch_val_541_453_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1309_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nfetch_val_453_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nfetch_val_453_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nfetch_val_453_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nfetch_val_453_Sample/ack
      -- 
    ack_1535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_541_453_buf_ack_0, ack => loadKernelChannel_CP_1309_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nfetch_val_453_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nfetch_val_453_Update/ack
      -- CP-element group 55: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nfetch_val_453_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_nfetch_val_453_Update/$exit
      -- 
    ack_1540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_541_453_buf_ack_1, ack => loadKernelChannel_CP_1309_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_my_fetch_454_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_my_fetch_454_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_my_fetch_454_sample_start__ps
      -- CP-element group 56: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_my_fetch_454_Sample/req
      -- 
    req_1552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(56), ack => my_fetch_414_454_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1309_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_my_fetch_454_update_start__ps
      -- CP-element group 57: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_my_fetch_454_Update/req
      -- CP-element group 57: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_my_fetch_454_update_start_
      -- CP-element group 57: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_my_fetch_454_Update/$entry
      -- 
    req_1557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(57), ack => my_fetch_414_454_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1309_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_my_fetch_454_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_my_fetch_454_sample_completed__ps
      -- CP-element group 58: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_my_fetch_454_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_my_fetch_454_Sample/ack
      -- 
    ack_1553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_414_454_buf_ack_0, ack => loadKernelChannel_CP_1309_elements(58)); -- 
    -- CP-element group 59:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_my_fetch_454_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_my_fetch_454_update_completed__ps
      -- CP-element group 59: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_my_fetch_454_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/R_my_fetch_454_Update/ack
      -- 
    ack_1558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_414_454_buf_ack_1, ack => loadKernelChannel_CP_1309_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	27 
    -- CP-element group 60: 	46 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe1_495_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe1_495_Sample/req
      -- CP-element group 60: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe1_495_Sample/$entry
      -- 
    req_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(60), ack => WPIPE_kernel_pipe1_495_inst_req_0); -- 
    loadKernelChannel_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(27) & loadKernelChannel_CP_1309_elements(46) & loadKernelChannel_CP_1309_elements(62);
      gj_loadKernelChannel_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	25 
    -- CP-element group 61: 	42 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe1_495_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe1_495_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe1_495_Sample/ack
      -- CP-element group 61: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe1_495_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe1_495_Update/req
      -- CP-element group 61: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe1_495_update_start_
      -- 
    ack_1568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_495_inst_ack_0, ack => loadKernelChannel_CP_1309_elements(61)); -- 
    req_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(61), ack => WPIPE_kernel_pipe1_495_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	93 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe1_495_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe1_495_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe1_495_Update/ack
      -- 
    ack_1573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_495_inst_ack_1, ack => loadKernelChannel_CP_1309_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	27 
    -- CP-element group 63: 	46 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe2_499_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe2_499_Sample/req
      -- CP-element group 63: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe2_499_Sample/$entry
      -- 
    req_1581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(63), ack => WPIPE_kernel_pipe2_499_inst_req_0); -- 
    loadKernelChannel_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(27) & loadKernelChannel_CP_1309_elements(46) & loadKernelChannel_CP_1309_elements(65);
      gj_loadKernelChannel_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	25 
    -- CP-element group 64: 	42 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe2_499_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe2_499_update_start_
      -- CP-element group 64: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe2_499_Update/req
      -- CP-element group 64: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe2_499_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe2_499_Sample/ack
      -- CP-element group 64: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe2_499_Update/$entry
      -- 
    ack_1582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_499_inst_ack_0, ack => loadKernelChannel_CP_1309_elements(64)); -- 
    req_1586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(64), ack => WPIPE_kernel_pipe2_499_inst_req_1); -- 
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	93 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	63 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe2_499_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe2_499_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe2_499_Update/ack
      -- 
    ack_1587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_499_inst_ack_1, ack => loadKernelChannel_CP_1309_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	27 
    -- CP-element group 66: 	46 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe3_503_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe3_503_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe3_503_Sample/req
      -- 
    req_1595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(66), ack => WPIPE_kernel_pipe3_503_inst_req_0); -- 
    loadKernelChannel_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(27) & loadKernelChannel_CP_1309_elements(46) & loadKernelChannel_CP_1309_elements(68);
      gj_loadKernelChannel_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	25 
    -- CP-element group 67: 	42 
    -- CP-element group 67:  members (6) 
      -- CP-element group 67: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe3_503_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe3_503_Update/req
      -- CP-element group 67: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe3_503_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe3_503_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe3_503_Sample/ack
      -- CP-element group 67: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe3_503_update_start_
      -- 
    ack_1596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe3_503_inst_ack_0, ack => loadKernelChannel_CP_1309_elements(67)); -- 
    req_1600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(67), ack => WPIPE_kernel_pipe3_503_inst_req_1); -- 
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	93 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	66 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe3_503_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe3_503_Update/ack
      -- CP-element group 68: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/WPIPE_kernel_pipe3_503_Update/$exit
      -- 
    ack_1601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe3_503_inst_ack_1, ack => loadKernelChannel_CP_1309_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	73 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	74 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	74 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/addr_of_520_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/addr_of_520_request/$entry
      -- CP-element group 69: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/addr_of_520_request/req
      -- 
    req_1641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(69), ack => addr_of_520_final_reg_req_0); -- 
    loadKernelChannel_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(73) & loadKernelChannel_CP_1309_elements(74);
      gj_loadKernelChannel_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	18 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	75 
    -- CP-element group 70: 	82 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	75 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/addr_of_520_update_start_
      -- CP-element group 70: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/addr_of_520_complete/$entry
      -- CP-element group 70: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/addr_of_520_complete/req
      -- 
    req_1646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(70), ack => addr_of_520_final_reg_req_1); -- 
    loadKernelChannel_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(18) & loadKernelChannel_CP_1309_elements(75) & loadKernelChannel_CP_1309_elements(82);
      gj_loadKernelChannel_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	18 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: 	74 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_final_index_sum_regn_update_start
      -- CP-element group 71: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_final_index_sum_regn_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_final_index_sum_regn_Update/req
      -- 
    req_1631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(71), ack => array_obj_ref_519_index_offset_req_1); -- 
    loadKernelChannel_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(18) & loadKernelChannel_CP_1309_elements(73) & loadKernelChannel_CP_1309_elements(74);
      gj_loadKernelChannel_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	27 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	93 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	25 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_final_index_sum_regn_sample_complete
      -- CP-element group 72: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_final_index_sum_regn_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_final_index_sum_regn_Sample/ack
      -- 
    ack_1627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_519_index_offset_ack_0, ack => loadKernelChannel_CP_1309_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	69 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (8) 
      -- CP-element group 73: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_offset_calculated
      -- CP-element group 73: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_final_index_sum_regn_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_final_index_sum_regn_Update/ack
      -- CP-element group 73: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/array_obj_ref_519_base_plus_offset/sum_rename_ack
      -- 
    ack_1632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_519_index_offset_ack_1, ack => loadKernelChannel_CP_1309_elements(73)); -- 
    -- CP-element group 74:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	69 
    -- CP-element group 74: successors 
    -- CP-element group 74: marked-successors 
    -- CP-element group 74: 	69 
    -- CP-element group 74: 	71 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/addr_of_520_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/addr_of_520_request/$exit
      -- CP-element group 74: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/addr_of_520_request/ack
      -- 
    ack_1642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_520_final_reg_ack_0, ack => loadKernelChannel_CP_1309_elements(74)); -- 
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	70 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	80 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	70 
    -- CP-element group 75:  members (19) 
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/addr_of_520_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_word_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/addr_of_520_complete/$exit
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/addr_of_520_complete/ack
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_base_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_root_address_calculated
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_base_address_resized
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_base_addr_resize/$entry
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_base_addr_resize/$exit
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_base_addr_resize/base_resize_req
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_base_addr_resize/base_resize_ack
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_base_plus_offset/$entry
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_base_plus_offset/$exit
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_base_plus_offset/sum_rename_req
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_base_plus_offset/sum_rename_ack
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_word_addrgen/$entry
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_word_addrgen/$exit
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_word_addrgen/root_register_req
      -- CP-element group 75: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_word_addrgen/root_register_ack
      -- 
    ack_1647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_520_final_reg_ack_1, ack => loadKernelChannel_CP_1309_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	27 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	78 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_524_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_524_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_524_Sample/req
      -- 
    req_1655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(76), ack => W_fn_486_delayed_7_0_522_inst_req_0); -- 
    loadKernelChannel_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(27) & loadKernelChannel_CP_1309_elements(78);
      gj_loadKernelChannel_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	79 
    -- CP-element group 77: 	82 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_524_update_start_
      -- CP-element group 77: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_524_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_524_Update/req
      -- 
    req_1660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(77), ack => W_fn_486_delayed_7_0_522_inst_req_1); -- 
    loadKernelChannel_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(79) & loadKernelChannel_CP_1309_elements(82);
      gj_loadKernelChannel_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	25 
    -- CP-element group 78: 	76 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_524_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_524_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_524_Sample/ack
      -- 
    ack_1656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_486_delayed_7_0_522_inst_ack_0, ack => loadKernelChannel_CP_1309_elements(78)); -- 
    -- CP-element group 79:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	77 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_524_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_524_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_524_Update/ack
      -- 
    ack_1661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_486_delayed_7_0_522_inst_ack_1, ack => loadKernelChannel_CP_1309_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	75 
    -- CP-element group 80: 	79 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Sample/word_access_start/$entry
      -- CP-element group 80: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Sample/word_access_start/word_0/$entry
      -- CP-element group 80: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Sample/word_access_start/word_0/rr
      -- 
    rr_1694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(80), ack => ptr_deref_528_load_0_req_0); -- 
    loadKernelChannel_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(75) & loadKernelChannel_CP_1309_elements(79) & loadKernelChannel_CP_1309_elements(82);
      gj_loadKernelChannel_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	21 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_update_start_
      -- CP-element group 81: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Update/word_access_complete/$entry
      -- CP-element group 81: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Update/word_access_complete/word_0/$entry
      -- CP-element group 81: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Update/word_access_complete/word_0/cr
      -- 
    cr_1705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(81), ack => ptr_deref_528_load_0_req_1); -- 
    loadKernelChannel_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(21) & loadKernelChannel_CP_1309_elements(83);
      gj_loadKernelChannel_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	70 
    -- CP-element group 82: 	77 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (5) 
      -- CP-element group 82: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Sample/word_access_start/$exit
      -- CP-element group 82: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Sample/word_access_start/word_0/$exit
      -- CP-element group 82: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Sample/word_access_start/word_0/ra
      -- 
    ra_1695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_528_load_0_ack_0, ack => loadKernelChannel_CP_1309_elements(82)); -- 
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	93 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	41 
    -- CP-element group 83: 	81 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Update/word_access_complete/$exit
      -- CP-element group 83: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Update/word_access_complete/word_0/$exit
      -- CP-element group 83: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Update/word_access_complete/word_0/ca
      -- CP-element group 83: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Update/ptr_deref_528_Merge/$entry
      -- CP-element group 83: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Update/ptr_deref_528_Merge/$exit
      -- CP-element group 83: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Update/ptr_deref_528_Merge/merge_req
      -- CP-element group 83: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/ptr_deref_528_Update/ptr_deref_528_Merge/merge_ack
      -- 
    ca_1706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_528_load_0_ack_1, ack => loadKernelChannel_CP_1309_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	27 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_532_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_532_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_532_Sample/req
      -- 
    req_1719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(84), ack => W_fn_492_delayed_13_0_530_inst_req_0); -- 
    loadKernelChannel_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(27) & loadKernelChannel_CP_1309_elements(86);
      gj_loadKernelChannel_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	21 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_532_update_start_
      -- CP-element group 85: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_532_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_532_Update/req
      -- 
    req_1724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(85), ack => W_fn_492_delayed_13_0_530_inst_req_1); -- 
    loadKernelChannel_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(21) & loadKernelChannel_CP_1309_elements(87);
      gj_loadKernelChannel_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	25 
    -- CP-element group 86: 	84 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_532_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_532_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_532_Sample/ack
      -- 
    ack_1720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_492_delayed_13_0_530_inst_ack_0, ack => loadKernelChannel_CP_1309_elements(86)); -- 
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	93 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	41 
    -- CP-element group 87: 	85 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_532_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_532_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_532_Update/ack
      -- 
    ack_1725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_492_delayed_13_0_530_inst_ack_1, ack => loadKernelChannel_CP_1309_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	46 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	90 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_535_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_535_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_535_Sample/req
      -- 
    req_1733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(88), ack => W_fetch_val_494_delayed_13_0_533_inst_req_0); -- 
    loadKernelChannel_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(46) & loadKernelChannel_CP_1309_elements(90);
      gj_loadKernelChannel_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	21 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_535_update_start_
      -- CP-element group 89: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_535_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_535_Update/req
      -- 
    req_1738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(89), ack => W_fetch_val_494_delayed_13_0_533_inst_req_1); -- 
    loadKernelChannel_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(21) & loadKernelChannel_CP_1309_elements(91);
      gj_loadKernelChannel_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	42 
    -- CP-element group 90: 	88 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_535_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_535_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_535_Sample/ack
      -- 
    ack_1734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_494_delayed_13_0_533_inst_ack_0, ack => loadKernelChannel_CP_1309_elements(90)); -- 
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	41 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_535_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_535_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/assign_stmt_535_Update/ack
      -- 
    ack_1739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_494_delayed_13_0_533_inst_ack_1, ack => loadKernelChannel_CP_1309_elements(91)); -- 
    -- CP-element group 92:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	18 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	19 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group loadKernelChannel_CP_1309_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => loadKernelChannel_CP_1309_elements(18), ack => loadKernelChannel_CP_1309_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  join  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	21 
    -- CP-element group 93: 	62 
    -- CP-element group 93: 	65 
    -- CP-element group 93: 	68 
    -- CP-element group 93: 	72 
    -- CP-element group 93: 	83 
    -- CP-element group 93: 	87 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	15 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_444/do_while_stmt_445/do_while_stmt_445_loop_body/$exit
      -- 
    loadKernelChannel_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1309_elements(91) & loadKernelChannel_CP_1309_elements(21) & loadKernelChannel_CP_1309_elements(62) & loadKernelChannel_CP_1309_elements(65) & loadKernelChannel_CP_1309_elements(68) & loadKernelChannel_CP_1309_elements(72) & loadKernelChannel_CP_1309_elements(83) & loadKernelChannel_CP_1309_elements(87);
      gj_loadKernelChannel_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	14 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_444/do_while_stmt_445/loop_exit/$exit
      -- CP-element group 94: 	 branch_block_stmt_444/do_while_stmt_445/loop_exit/ack
      -- 
    ack_1744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_445_branch_ack_0, ack => loadKernelChannel_CP_1309_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	14 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_444/do_while_stmt_445/loop_taken/$exit
      -- CP-element group 95: 	 branch_block_stmt_444/do_while_stmt_445/loop_taken/ack
      -- 
    ack_1748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_445_branch_ack_1, ack => loadKernelChannel_CP_1309_elements(95)); -- 
    -- CP-element group 96:  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	12 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	10 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_444/do_while_stmt_445/$exit
      -- 
    loadKernelChannel_CP_1309_elements(96) <= loadKernelChannel_CP_1309_elements(12);
    -- CP-element group 97:  transition  input  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	10 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (6) 
      -- CP-element group 97: 	 assign_stmt_551/WPIPE_size_pipe_549_sample_completed_
      -- CP-element group 97: 	 assign_stmt_551/WPIPE_size_pipe_549_update_start_
      -- CP-element group 97: 	 assign_stmt_551/WPIPE_size_pipe_549_Sample/$exit
      -- CP-element group 97: 	 assign_stmt_551/WPIPE_size_pipe_549_Sample/ack
      -- CP-element group 97: 	 assign_stmt_551/WPIPE_size_pipe_549_Update/$entry
      -- CP-element group 97: 	 assign_stmt_551/WPIPE_size_pipe_549_Update/req
      -- 
    ack_1761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_549_inst_ack_0, ack => loadKernelChannel_CP_1309_elements(97)); -- 
    req_1765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1309_elements(97), ack => WPIPE_size_pipe_549_inst_req_1); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (5) 
      -- CP-element group 98: 	 $exit
      -- CP-element group 98: 	 assign_stmt_551/$exit
      -- CP-element group 98: 	 assign_stmt_551/WPIPE_size_pipe_549_update_completed_
      -- CP-element group 98: 	 assign_stmt_551/WPIPE_size_pipe_549_Update/$exit
      -- CP-element group 98: 	 assign_stmt_551/WPIPE_size_pipe_549_Update/ack
      -- 
    ack_1766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_549_inst_ack_1, ack => loadKernelChannel_CP_1309_elements(98)); -- 
    loadKernelChannel_do_while_stmt_445_terminator_1749: loop_terminator -- 
      generic map (name => " loadKernelChannel_do_while_stmt_445_terminator_1749", max_iterations_in_flight =>15) 
      port map(loop_body_exit => loadKernelChannel_CP_1309_elements(15),loop_continue => loadKernelChannel_CP_1309_elements(95),loop_terminate => loadKernelChannel_CP_1309_elements(94),loop_back => loadKernelChannel_CP_1309_elements(13),loop_exit => loadKernelChannel_CP_1309_elements(12),clk => clk, reset => reset); -- 
    phi_stmt_447_phi_seq_1505_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_1309_elements(30);
      loadKernelChannel_CP_1309_elements(33)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_1309_elements(35);
      loadKernelChannel_CP_1309_elements(34)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_1309_elements(36);
      loadKernelChannel_CP_1309_elements(31) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_1309_elements(28);
      loadKernelChannel_CP_1309_elements(37)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_1309_elements(39);
      loadKernelChannel_CP_1309_elements(38)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_1309_elements(40);
      loadKernelChannel_CP_1309_elements(29) <= phi_mux_reqs(1);
      phi_stmt_447_phi_seq_1505 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_447_phi_seq_1505") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_1309_elements(20), 
          phi_sample_ack => loadKernelChannel_CP_1309_elements(26), 
          phi_update_req => loadKernelChannel_CP_1309_elements(22), 
          phi_update_ack => loadKernelChannel_CP_1309_elements(27), 
          phi_mux_ack => loadKernelChannel_CP_1309_elements(32), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_451_phi_seq_1559_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_1309_elements(47);
      loadKernelChannel_CP_1309_elements(52)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_1309_elements(54);
      loadKernelChannel_CP_1309_elements(53)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_1309_elements(55);
      loadKernelChannel_CP_1309_elements(48) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_1309_elements(49);
      loadKernelChannel_CP_1309_elements(56)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_1309_elements(58);
      loadKernelChannel_CP_1309_elements(57)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_1309_elements(59);
      loadKernelChannel_CP_1309_elements(50) <= phi_mux_reqs(1);
      phi_stmt_451_phi_seq_1559 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_451_phi_seq_1559") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_1309_elements(43), 
          phi_sample_ack => loadKernelChannel_CP_1309_elements(44), 
          phi_update_req => loadKernelChannel_CP_1309_elements(45), 
          phi_update_ack => loadKernelChannel_CP_1309_elements(46), 
          phi_mux_ack => loadKernelChannel_CP_1309_elements(51), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1447_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= loadKernelChannel_CP_1309_elements(16);
        preds(1)  <= loadKernelChannel_CP_1309_elements(17);
        entry_tmerge_1447 : transition_merge -- 
          generic map(name => " entry_tmerge_1447")
          port map (preds => preds, symbol_out => loadKernelChannel_CP_1309_elements(18));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u64_u64_460_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_509_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_473_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_518_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_518_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_518_wire : std_logic_vector(63 downto 0);
    signal NOT_u1_u1_483_wire : std_logic_vector(0 downto 0);
    signal R_sh_start_407_resized : std_logic_vector(13 downto 0);
    signal R_sh_start_407_scaled : std_logic_vector(13 downto 0);
    signal SHL_u16_u16_396_wire : std_logic_vector(15 downto 0);
    signal SHL_u16_u16_425_wire : std_logic_vector(15 downto 0);
    signal SUB_u64_u64_461_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_546_wire : std_logic_vector(63 downto 0);
    signal ULT_u64_u1_486_wire : std_logic_vector(0 downto 0);
    signal ULT_u64_u1_547_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_408_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_408_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_408_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_408_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_408_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_408_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_519_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_519_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_519_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_519_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_519_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_519_root_address : std_logic_vector(13 downto 0);
    signal ea1_420 : std_logic_vector(63 downto 0);
    signal ea2_428 : std_logic_vector(63 downto 0);
    signal ea3_434 : std_logic_vector(63 downto 0);
    signal fetch_addr_410 : std_logic_vector(31 downto 0);
    signal fetch_addr_521 : std_logic_vector(31 downto 0);
    signal fetch_val_451 : std_logic_vector(63 downto 0);
    signal fetch_val_494_delayed_13_0_535 : std_logic_vector(63 downto 0);
    signal first_fill_439 : std_logic_vector(0 downto 0);
    signal fn_486_delayed_7_0_524 : std_logic_vector(0 downto 0);
    signal fn_492_delayed_13_0_532 : std_logic_vector(0 downto 0);
    signal fn_512 : std_logic_vector(0 downto 0);
    signal fv_529 : std_logic_vector(63 downto 0);
    signal konst_395_wire_constant : std_logic_vector(15 downto 0);
    signal konst_401_wire_constant : std_logic_vector(63 downto 0);
    signal konst_424_wire_constant : std_logic_vector(15 downto 0);
    signal konst_437_wire_constant : std_logic_vector(63 downto 0);
    signal konst_457_wire_constant : std_logic_vector(63 downto 0);
    signal konst_459_wire_constant : std_logic_vector(63 downto 0);
    signal konst_462_wire_constant : std_logic_vector(63 downto 0);
    signal konst_467_wire_constant : std_logic_vector(63 downto 0);
    signal konst_508_wire_constant : std_logic_vector(63 downto 0);
    signal konst_510_wire_constant : std_logic_vector(63 downto 0);
    signal konst_517_wire_constant : std_logic_vector(63 downto 0);
    signal konst_545_wire_constant : std_logic_vector(63 downto 0);
    signal my_fetch_414 : std_logic_vector(63 downto 0);
    signal my_fetch_414_454_buffered : std_logic_vector(63 downto 0);
    signal my_num1_464 : std_logic_vector(63 downto 0);
    signal mycount_447 : std_logic_vector(63 downto 0);
    signal nfetch_val_541 : std_logic_vector(63 downto 0);
    signal nfetch_val_541_453_buffered : std_logic_vector(63 downto 0);
    signal nmycount_469 : std_logic_vector(63 downto 0);
    signal nmycount_469_450_buffered : std_logic_vector(63 downto 0);
    signal ptr_deref_413_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_413_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_413_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_413_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_413_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_528_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_528_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_528_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_528_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_528_word_offset_0 : std_logic_vector(13 downto 0);
    signal row_size_398 : std_logic_vector(15 downto 0);
    signal send_to_1_480 : std_logic_vector(0 downto 0);
    signal send_to_2_488 : std_logic_vector(0 downto 0);
    signal send_to_3_493 : std_logic_vector(0 downto 0);
    signal sh_start_403 : std_logic_vector(63 downto 0);
    signal start_add_449_buffered : std_logic_vector(63 downto 0);
    signal start_next_443 : std_logic_vector(7 downto 0);
    signal type_cast_418_wire : std_logic_vector(63 downto 0);
    signal type_cast_426_wire : std_logic_vector(63 downto 0);
    signal type_cast_432_wire : std_logic_vector(63 downto 0);
    signal var_val_475 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_408_constant_part_of_offset <= "00000000000000";
    array_obj_ref_408_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_408_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_408_resized_base_address <= "00000000000000";
    array_obj_ref_519_constant_part_of_offset <= "00000000000000";
    array_obj_ref_519_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_519_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_519_resized_base_address <= "00000000000000";
    konst_395_wire_constant <= "0000000000000001";
    konst_401_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_424_wire_constant <= "0000000000000001";
    konst_437_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_457_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_459_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_462_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_467_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_508_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_510_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_517_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_545_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    ptr_deref_413_word_offset_0 <= "00000000000000";
    ptr_deref_528_word_offset_0 <= "00000000000000";
    phi_stmt_447: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= start_add_449_buffered & nmycount_469_450_buffered;
      req <= phi_stmt_447_req_0 & phi_stmt_447_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_447",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_447_ack_0,
          idata => idata,
          odata => mycount_447,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_447
    phi_stmt_451: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nfetch_val_541_453_buffered & my_fetch_414_454_buffered;
      req <= phi_stmt_451_req_0 & phi_stmt_451_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_451",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_451_ack_0,
          idata => idata,
          odata => fetch_val_451,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_451
    -- flow-through select operator MUX_540_inst
    nfetch_val_541 <= fv_529 when (fn_492_delayed_13_0_532(0) /=  '0') else fetch_val_494_delayed_13_0_535;
    W_fetch_val_494_delayed_13_0_533_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val_494_delayed_13_0_533_inst_req_0;
      W_fetch_val_494_delayed_13_0_533_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val_494_delayed_13_0_533_inst_req_1;
      W_fetch_val_494_delayed_13_0_533_inst_ack_1<= rack(0);
      W_fetch_val_494_delayed_13_0_533_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val_494_delayed_13_0_533_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val_451,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val_494_delayed_13_0_535,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_486_delayed_7_0_522_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_486_delayed_7_0_522_inst_req_0;
      W_fn_486_delayed_7_0_522_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_486_delayed_7_0_522_inst_req_1;
      W_fn_486_delayed_7_0_522_inst_ack_1<= rack(0);
      W_fn_486_delayed_7_0_522_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_486_delayed_7_0_522_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_512,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_486_delayed_7_0_524,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_492_delayed_13_0_530_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_492_delayed_13_0_530_inst_req_0;
      W_fn_492_delayed_13_0_530_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_492_delayed_13_0_530_inst_req_1;
      W_fn_492_delayed_13_0_530_inst_ack_1<= rack(0);
      W_fn_492_delayed_13_0_530_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_492_delayed_13_0_530_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_512,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_492_delayed_13_0_532,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_409_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_409_final_reg_req_0;
      addr_of_409_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_409_final_reg_req_1;
      addr_of_409_final_reg_ack_1<= rack(0);
      addr_of_409_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_409_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_408_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_410,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_520_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_520_final_reg_req_0;
      addr_of_520_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_520_final_reg_req_1;
      addr_of_520_final_reg_ack_1<= rack(0);
      addr_of_520_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_520_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_519_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_521,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch_414_454_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch_414_454_buf_req_0;
      my_fetch_414_454_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch_414_454_buf_req_1;
      my_fetch_414_454_buf_ack_1<= rack(0);
      my_fetch_414_454_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch_414_454_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch_414,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch_414_454_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nfetch_val_541_453_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nfetch_val_541_453_buf_req_0;
      nfetch_val_541_453_buf_ack_0<= wack(0);
      rreq(0) <= nfetch_val_541_453_buf_req_1;
      nfetch_val_541_453_buf_ack_1<= rack(0);
      nfetch_val_541_453_buf : InterlockBuffer generic map ( -- 
        name => "nfetch_val_541_453_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nfetch_val_541,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nfetch_val_541_453_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_469_450_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_469_450_buf_req_0;
      nmycount_469_450_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_469_450_buf_req_1;
      nmycount_469_450_buf_ack_1<= rack(0);
      nmycount_469_450_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_469_450_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_469,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_469_450_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    start_add_449_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= start_add_449_buf_req_0;
      start_add_449_buf_ack_0<= wack(0);
      rreq(0) <= start_add_449_buf_req_1;
      start_add_449_buf_ack_1<= rack(0);
      start_add_449_buf : InterlockBuffer generic map ( -- 
        name => "start_add_449_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => start_add_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => start_add_449_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_418_inst
    process(row_size_398) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := row_size_398(15 downto 0);
      type_cast_418_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_426_inst
    process(SHL_u16_u16_425_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := SHL_u16_u16_425_wire(15 downto 0);
      type_cast_426_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_432_inst
    process(row_size_398) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := row_size_398(15 downto 0);
      type_cast_432_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_474_inst
    process(LSHR_u64_u64_473_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_473_wire(15 downto 0);
      var_val_475 <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_408_index_1_rename
    process(R_sh_start_407_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_sh_start_407_resized;
      ov(13 downto 0) := iv;
      R_sh_start_407_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_408_index_1_resize
    process(sh_start_403) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := sh_start_403;
      ov := iv(13 downto 0);
      R_sh_start_407_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_408_root_address_inst
    process(array_obj_ref_408_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_408_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_408_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_519_index_1_rename
    process(LSHR_u64_u64_518_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_518_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_518_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_519_index_1_resize
    process(LSHR_u64_u64_518_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_518_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_518_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_519_root_address_inst
    process(array_obj_ref_519_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_519_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_519_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_413_addr_0
    process(ptr_deref_413_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_413_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_413_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_413_base_resize
    process(fetch_addr_410) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_410;
      ov := iv(13 downto 0);
      ptr_deref_413_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_413_gather_scatter
    process(ptr_deref_413_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_413_data_0;
      ov(63 downto 0) := iv;
      my_fetch_414 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_413_root_address_inst
    process(ptr_deref_413_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_413_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_413_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_528_addr_0
    process(ptr_deref_528_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_528_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_528_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_528_base_resize
    process(fetch_addr_521) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_521;
      ov := iv(13 downto 0);
      ptr_deref_528_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_528_gather_scatter
    process(ptr_deref_528_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_528_data_0;
      ov(63 downto 0) := iv;
      fv_529 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_528_root_address_inst
    process(ptr_deref_528_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_528_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_528_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_445_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u64_u1_547_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_445_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_445_branch_req_0,
          ack0 => do_while_stmt_445_branch_ack_0,
          ack1 => do_while_stmt_445_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_397_inst
    process(num_chl_buffer, SHL_u16_u16_396_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_chl_buffer, SHL_u16_u16_396_wire, tmp_var);
      row_size_398 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_419_inst
    process(start_add_buffer, type_cast_418_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(start_add_buffer, type_cast_418_wire, tmp_var);
      ea1_420 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_427_inst
    process(start_add_buffer, type_cast_426_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(start_add_buffer, type_cast_426_wire, tmp_var);
      ea2_428 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_433_inst
    process(ea2_428, type_cast_432_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ea2_428, type_cast_432_wire, tmp_var);
      ea3_434 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_468_inst
    process(mycount_447) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_447, konst_467_wire_constant, tmp_var);
      nmycount_469 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_487_inst
    process(NOT_u1_u1_483_wire, ULT_u64_u1_486_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_483_wire, ULT_u64_u1_486_wire, tmp_var);
      send_to_2_488 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_460_inst
    process(mycount_447) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mycount_447, konst_459_wire_constant, tmp_var);
      AND_u64_u64_460_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_509_inst
    process(nmycount_469) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(nmycount_469, konst_508_wire_constant, tmp_var);
      AND_u64_u64_509_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_438_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(start_add_buffer, konst_437_wire_constant, tmp_var);
      first_fill_439 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_511_inst
    process(AND_u64_u64_509_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(AND_u64_u64_509_wire, konst_510_wire_constant, tmp_var);
      fn_512 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_402_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(start_add_buffer, konst_401_wire_constant, tmp_var);
      sh_start_403 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_473_inst
    process(fetch_val_451, my_num1_464) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val_451, my_num1_464, tmp_var);
      LSHR_u64_u64_473_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_518_inst
    process(nmycount_469) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(nmycount_469, konst_517_wire_constant, tmp_var);
      LSHR_u64_u64_518_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_483_inst
    process(send_to_1_480) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", send_to_1_480, tmp_var);
      NOT_u1_u1_483_wire <= tmp_var; -- 
    end process;
    -- binary operator SHL_u16_u16_396_inst
    process(num_chl_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(num_chl_buffer, konst_395_wire_constant, tmp_var);
      SHL_u16_u16_396_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_425_inst
    process(row_size_398) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(row_size_398, konst_424_wire_constant, tmp_var);
      SHL_u16_u16_425_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_463_inst
    process(SUB_u64_u64_461_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_461_wire, konst_462_wire_constant, tmp_var);
      my_num1_464 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_461_inst
    process(konst_457_wire_constant, AND_u64_u64_460_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_457_wire_constant, AND_u64_u64_460_wire, tmp_var);
      SUB_u64_u64_461_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_546_inst
    process(ea3_434) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(ea3_434, konst_545_wire_constant, tmp_var);
      SUB_u64_u64_546_wire <= tmp_var; --
    end process;
    -- binary operator UGE_u64_u1_492_inst
    process(mycount_447, ea2_428) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(mycount_447, ea2_428, tmp_var);
      send_to_3_493 <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_479_inst
    process(mycount_447, ea1_420) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_447, ea1_420, tmp_var);
      send_to_1_480 <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_486_inst
    process(mycount_447, ea2_428) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_447, ea2_428, tmp_var);
      ULT_u64_u1_486_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_547_inst
    process(mycount_447, SUB_u64_u64_546_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_447, SUB_u64_u64_546_wire, tmp_var);
      ULT_u64_u1_547_wire <= tmp_var; --
    end process;
    -- shared split operator group (23) : array_obj_ref_408_index_offset 
    ApIntAdd_group_23: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_sh_start_407_scaled;
      array_obj_ref_408_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_408_index_offset_req_0;
      array_obj_ref_408_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_408_index_offset_req_1;
      array_obj_ref_408_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_23_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_23_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_23",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : array_obj_ref_519_index_offset 
    ApIntAdd_group_24: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_518_scaled;
      array_obj_ref_519_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_519_index_offset_req_0;
      array_obj_ref_519_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_519_index_offset_req_1;
      array_obj_ref_519_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_24_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_24_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_24",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared load operator group (0) : ptr_deref_528_load_0 ptr_deref_413_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 6);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_528_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_413_load_0_req_0;
      ptr_deref_528_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_413_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_528_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_413_load_0_req_1;
      ptr_deref_528_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_413_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <= fn_486_delayed_7_0_524(0);
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_528_word_address_0 & ptr_deref_413_word_address_0;
      ptr_deref_528_data_0 <= data_out(127 downto 64);
      ptr_deref_413_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_input_done_pipe_442_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_done_pipe_442_inst_req_0;
      RPIPE_input_done_pipe_442_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_done_pipe_442_inst_req_1;
      RPIPE_input_done_pipe_442_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not first_fill_439(0);
      start_next_443 <= data_out(7 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_kernel_pipe1_495_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_495_inst_req_0;
      WPIPE_kernel_pipe1_495_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_495_inst_req_1;
      WPIPE_kernel_pipe1_495_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_480(0);
      data_in <= var_val_475;
      kernel_pipe1_write_0_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_kernel_pipe2_499_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe2_499_inst_req_0;
      WPIPE_kernel_pipe2_499_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe2_499_inst_req_1;
      WPIPE_kernel_pipe2_499_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_488(0);
      data_in <= var_val_475;
      kernel_pipe2_write_1_gI: SplitGuardInterface generic map(name => "kernel_pipe2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe2_write_1: OutputPortRevised -- 
        generic map ( name => "kernel_pipe2", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe2_pipe_write_req(0),
          oack => kernel_pipe2_pipe_write_ack(0),
          odata => kernel_pipe2_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_kernel_pipe3_503_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe3_503_inst_req_0;
      WPIPE_kernel_pipe3_503_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe3_503_inst_req_1;
      WPIPE_kernel_pipe3_503_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_493(0);
      data_in <= var_val_475;
      kernel_pipe3_write_2_gI: SplitGuardInterface generic map(name => "kernel_pipe3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe3_write_2: OutputPortRevised -- 
        generic map ( name => "kernel_pipe3", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe3_pipe_write_req(0),
          oack => kernel_pipe3_pipe_write_ack(0),
          odata => kernel_pipe3_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_size_pipe_549_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_size_pipe_549_inst_req_0;
      WPIPE_size_pipe_549_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_size_pipe_549_inst_req_1;
      WPIPE_size_pipe_549_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= num_chl_buffer;
      size_pipe_write_3_gI: SplitGuardInterface generic map(name => "size_pipe_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      size_pipe_write_3: OutputPortRevised -- 
        generic map ( name => "size_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => size_pipe_pipe_write_req(0),
          oack => size_pipe_pipe_write_ack(0),
          odata => size_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end loadKernelChannel_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_1275_start: Boolean;
  signal timer_CP_1275_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_req_381_inst_req_0 : boolean;
  signal WPIPE_timer_req_381_inst_ack_0 : boolean;
  signal WPIPE_timer_req_381_inst_req_1 : boolean;
  signal WPIPE_timer_req_381_inst_ack_1 : boolean;
  signal RPIPE_timer_resp_386_inst_req_0 : boolean;
  signal RPIPE_timer_resp_386_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_386_inst_req_1 : boolean;
  signal RPIPE_timer_resp_386_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_1275_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_1275_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_1275_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_1275_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_1275: Block -- control-path 
    signal timer_CP_1275_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_1275_elements(0) <= timer_CP_1275_start;
    timer_CP_1275_symbol <= timer_CP_1275_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_384_to_assign_stmt_387/$entry
      -- CP-element group 0: 	 assign_stmt_384_to_assign_stmt_387/WPIPE_timer_req_381_sample_start_
      -- CP-element group 0: 	 assign_stmt_384_to_assign_stmt_387/WPIPE_timer_req_381_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_384_to_assign_stmt_387/WPIPE_timer_req_381_Sample/req
      -- CP-element group 0: 	 assign_stmt_384_to_assign_stmt_387/RPIPE_timer_resp_386_sample_start_
      -- CP-element group 0: 	 assign_stmt_384_to_assign_stmt_387/RPIPE_timer_resp_386_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_384_to_assign_stmt_387/RPIPE_timer_resp_386_Sample/rr
      -- 
    req_1288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1275_elements(0), ack => WPIPE_timer_req_381_inst_req_0); -- 
    rr_1302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1275_elements(0), ack => RPIPE_timer_resp_386_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_384_to_assign_stmt_387/WPIPE_timer_req_381_sample_completed_
      -- CP-element group 1: 	 assign_stmt_384_to_assign_stmt_387/WPIPE_timer_req_381_update_start_
      -- CP-element group 1: 	 assign_stmt_384_to_assign_stmt_387/WPIPE_timer_req_381_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_384_to_assign_stmt_387/WPIPE_timer_req_381_Sample/ack
      -- CP-element group 1: 	 assign_stmt_384_to_assign_stmt_387/WPIPE_timer_req_381_Update/$entry
      -- CP-element group 1: 	 assign_stmt_384_to_assign_stmt_387/WPIPE_timer_req_381_Update/req
      -- 
    ack_1289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_381_inst_ack_0, ack => timer_CP_1275_elements(1)); -- 
    req_1293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1275_elements(1), ack => WPIPE_timer_req_381_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_384_to_assign_stmt_387/WPIPE_timer_req_381_update_completed_
      -- CP-element group 2: 	 assign_stmt_384_to_assign_stmt_387/WPIPE_timer_req_381_Update/$exit
      -- CP-element group 2: 	 assign_stmt_384_to_assign_stmt_387/WPIPE_timer_req_381_Update/ack
      -- 
    ack_1294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_381_inst_ack_1, ack => timer_CP_1275_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_384_to_assign_stmt_387/RPIPE_timer_resp_386_sample_completed_
      -- CP-element group 3: 	 assign_stmt_384_to_assign_stmt_387/RPIPE_timer_resp_386_update_start_
      -- CP-element group 3: 	 assign_stmt_384_to_assign_stmt_387/RPIPE_timer_resp_386_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_384_to_assign_stmt_387/RPIPE_timer_resp_386_Sample/ra
      -- CP-element group 3: 	 assign_stmt_384_to_assign_stmt_387/RPIPE_timer_resp_386_Update/$entry
      -- CP-element group 3: 	 assign_stmt_384_to_assign_stmt_387/RPIPE_timer_resp_386_Update/cr
      -- 
    ra_1303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_386_inst_ack_0, ack => timer_CP_1275_elements(3)); -- 
    cr_1307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1275_elements(3), ack => RPIPE_timer_resp_386_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_384_to_assign_stmt_387/RPIPE_timer_resp_386_update_completed_
      -- CP-element group 4: 	 assign_stmt_384_to_assign_stmt_387/RPIPE_timer_resp_386_Update/$exit
      -- CP-element group 4: 	 assign_stmt_384_to_assign_stmt_387/RPIPE_timer_resp_386_Update/ca
      -- 
    ca_1308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_386_inst_ack_1, ack => timer_CP_1275_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_384_to_assign_stmt_387/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_1275_elements(2) & timer_CP_1275_elements(4);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_1275_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_383_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_383_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_386_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_386_inst_req_0;
      RPIPE_timer_resp_386_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_386_inst_req_1;
      RPIPE_timer_resp_386_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_381_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_381_inst_req_0;
      WPIPE_timer_req_381_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_381_inst_req_1;
      WPIPE_timer_req_381_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_383_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_5950_start: Boolean;
  signal timerDaemon_CP_5950_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_resp_2450_inst_ack_0 : boolean;
  signal WPIPE_timer_resp_2450_inst_req_0 : boolean;
  signal phi_stmt_2435_req_1 : boolean;
  signal WPIPE_timer_resp_2450_inst_req_1 : boolean;
  signal WPIPE_timer_resp_2450_inst_ack_1 : boolean;
  signal phi_stmt_2435_req_0 : boolean;
  signal nCOUNTER_2448_2439_buf_req_0 : boolean;
  signal phi_stmt_2435_ack_0 : boolean;
  signal do_while_stmt_2433_branch_ack_0 : boolean;
  signal RPIPE_timer_req_2442_inst_ack_1 : boolean;
  signal RPIPE_timer_req_2442_inst_req_1 : boolean;
  signal RPIPE_timer_req_2442_inst_ack_0 : boolean;
  signal RPIPE_timer_req_2442_inst_req_0 : boolean;
  signal do_while_stmt_2433_branch_ack_1 : boolean;
  signal nCOUNTER_2448_2439_buf_ack_1 : boolean;
  signal do_while_stmt_2433_branch_req_0 : boolean;
  signal nCOUNTER_2448_2439_buf_req_1 : boolean;
  signal nCOUNTER_2448_2439_buf_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_5950_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_5950_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_5950_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_5950_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_5950: Block -- control-path 
    signal timerDaemon_CP_5950_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_5950_elements(0) <= timerDaemon_CP_5950_start;
    timerDaemon_CP_5950_symbol <= timerDaemon_CP_5950_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2432/$entry
      -- CP-element group 0: 	 branch_block_stmt_2432/do_while_stmt_2433__entry__
      -- CP-element group 0: 	 branch_block_stmt_2432/branch_block_stmt_2432__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_2432/do_while_stmt_2433__exit__
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_2432/$exit
      -- CP-element group 1: 	 branch_block_stmt_2432/branch_block_stmt_2432__exit__
      -- 
    timerDaemon_CP_5950_elements(1) <= timerDaemon_CP_5950_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433__entry__
      -- CP-element group 2: 	 branch_block_stmt_2432/do_while_stmt_2433/$entry
      -- 
    timerDaemon_CP_5950_elements(2) <= timerDaemon_CP_5950_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433__exit__
      -- 
    -- Element group timerDaemon_CP_5950_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_2432/do_while_stmt_2433/loop_back
      -- 
    -- Element group timerDaemon_CP_5950_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: 	43 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2432/do_while_stmt_2433/condition_done
      -- CP-element group 5: 	 branch_block_stmt_2432/do_while_stmt_2433/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_2432/do_while_stmt_2433/loop_taken/$entry
      -- 
    timerDaemon_CP_5950_elements(5) <= timerDaemon_CP_5950_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_2432/do_while_stmt_2433/loop_body_done
      -- 
    timerDaemon_CP_5950_elements(6) <= timerDaemon_CP_5950_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_5950_elements(7) <= timerDaemon_CP_5950_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_5950_elements(8) <= timerDaemon_CP_5950_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	40 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2440_sample_start_
      -- 
    -- Element group timerDaemon_CP_5950_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	40 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/condition_evaluated
      -- 
    condition_evaluated_5974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_5974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5950_elements(10), ack => do_while_stmt_2433_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5950_elements(14) & timerDaemon_CP_5950_elements(40);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5950_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2435_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/aggregated_phi_sample_req
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_5950_elements(9) & timerDaemon_CP_5950_elements(15) & timerDaemon_CP_5950_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5950_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	35 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2435_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2440_sample_completed_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5950_elements(17) & timerDaemon_CP_5950_elements(35);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5950_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2435_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/aggregated_phi_update_req
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5950_elements(16) & timerDaemon_CP_5950_elements(32);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5950_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	36 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5950_elements(18) & timerDaemon_CP_5950_elements(36);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5950_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2435_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5950_elements(9) & timerDaemon_CP_5950_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5950_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2435_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5950_elements(9) & timerDaemon_CP_5950_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5950_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2435_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_5950_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	37 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2435_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2435_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_5950_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2435_loopback_trigger
      -- 
    timerDaemon_CP_5950_elements(19) <= timerDaemon_CP_5950_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2435_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2435_loopback_sample_req_ps
      -- 
    phi_stmt_2435_loopback_sample_req_5989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2435_loopback_sample_req_5989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5950_elements(20), ack => phi_stmt_2435_req_1); -- 
    -- Element group timerDaemon_CP_5950_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2435_entry_trigger
      -- 
    timerDaemon_CP_5950_elements(21) <= timerDaemon_CP_5950_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2435_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2435_entry_sample_req_ps
      -- 
    phi_stmt_2435_entry_sample_req_5992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2435_entry_sample_req_5992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5950_elements(22), ack => phi_stmt_2435_req_0); -- 
    -- Element group timerDaemon_CP_5950_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2435_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2435_phi_mux_ack_ps
      -- 
    phi_stmt_2435_phi_mux_ack_5995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2435_ack_0, ack => timerDaemon_CP_5950_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/type_cast_2438_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/type_cast_2438_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/type_cast_2438_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/type_cast_2438_sample_completed_
      -- 
    -- Element group timerDaemon_CP_5950_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/type_cast_2438_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/type_cast_2438_update_start_
      -- 
    -- Element group timerDaemon_CP_5950_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/type_cast_2438_update_completed__ps
      -- 
    timerDaemon_CP_5950_elements(26) <= timerDaemon_CP_5950_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/type_cast_2438_update_completed_
      -- 
    -- Element group timerDaemon_CP_5950_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => timerDaemon_CP_5950_elements(25), ack => timerDaemon_CP_5950_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/R_nCOUNTER_2439_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/R_nCOUNTER_2439_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/R_nCOUNTER_2439_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/R_nCOUNTER_2439_sample_start__ps
      -- 
    req_6016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5950_elements(28), ack => nCOUNTER_2448_2439_buf_req_0); -- 
    -- Element group timerDaemon_CP_5950_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/R_nCOUNTER_2439_update_start_
      -- CP-element group 29: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/R_nCOUNTER_2439_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/R_nCOUNTER_2439_Update/req
      -- CP-element group 29: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/R_nCOUNTER_2439_Update/$entry
      -- 
    req_6021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5950_elements(29), ack => nCOUNTER_2448_2439_buf_req_1); -- 
    -- Element group timerDaemon_CP_5950_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/R_nCOUNTER_2439_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/R_nCOUNTER_2439_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/R_nCOUNTER_2439_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/R_nCOUNTER_2439_Sample/ack
      -- 
    ack_6017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_2448_2439_buf_ack_0, ack => timerDaemon_CP_5950_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/R_nCOUNTER_2439_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/R_nCOUNTER_2439_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/R_nCOUNTER_2439_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/R_nCOUNTER_2439_Update/$exit
      -- 
    ack_6022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_2448_2439_buf_ack_1, ack => timerDaemon_CP_5950_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2440_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5950_elements(9) & timerDaemon_CP_5950_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5950_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/RPIPE_timer_req_2442_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/RPIPE_timer_req_2442_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/RPIPE_timer_req_2442_sample_start_
      -- 
    rr_6035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5950_elements(33), ack => RPIPE_timer_req_2442_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5950_elements(11) & timerDaemon_CP_5950_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5950_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	13 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/RPIPE_timer_req_2442_Update/cr
      -- CP-element group 34: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/RPIPE_timer_req_2442_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/RPIPE_timer_req_2442_update_start_
      -- 
    cr_6040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5950_elements(34), ack => RPIPE_timer_req_2442_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5950_elements(13) & timerDaemon_CP_5950_elements(35);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5950_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/RPIPE_timer_req_2442_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/RPIPE_timer_req_2442_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/RPIPE_timer_req_2442_sample_completed_
      -- 
    ra_6036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_2442_inst_ack_0, ack => timerDaemon_CP_5950_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: 	37 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/RPIPE_timer_req_2442_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/RPIPE_timer_req_2442_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/RPIPE_timer_req_2442_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/phi_stmt_2440_update_completed_
      -- 
    ca_6041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_2442_inst_ack_1, ack => timerDaemon_CP_5950_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	18 
    -- CP-element group 37: 	36 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/WPIPE_timer_resp_2450_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/WPIPE_timer_resp_2450_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/WPIPE_timer_resp_2450_sample_start_
      -- 
    req_6049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5950_elements(37), ack => WPIPE_timer_resp_2450_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_5950_elements(18) & timerDaemon_CP_5950_elements(36) & timerDaemon_CP_5950_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5950_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	16 
    -- CP-element group 38: 	32 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/WPIPE_timer_resp_2450_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/WPIPE_timer_resp_2450_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/WPIPE_timer_resp_2450_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/WPIPE_timer_resp_2450_Update/req
      -- CP-element group 38: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/WPIPE_timer_resp_2450_update_start_
      -- CP-element group 38: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/WPIPE_timer_resp_2450_sample_completed_
      -- 
    ack_6050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_2450_inst_ack_0, ack => timerDaemon_CP_5950_elements(38)); -- 
    req_6054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5950_elements(38), ack => WPIPE_timer_resp_2450_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/WPIPE_timer_resp_2450_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/WPIPE_timer_resp_2450_Update/ack
      -- CP-element group 39: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/WPIPE_timer_resp_2450_update_completed_
      -- 
    ack_6055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_2450_inst_ack_1, ack => timerDaemon_CP_5950_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_5950_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_5950_elements(9), ack => timerDaemon_CP_5950_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	12 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_2432/do_while_stmt_2433/do_while_stmt_2433_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5950_elements(12) & timerDaemon_CP_5950_elements(39);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5950_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_2432/do_while_stmt_2433/loop_exit/$exit
      -- CP-element group 42: 	 branch_block_stmt_2432/do_while_stmt_2433/loop_exit/ack
      -- 
    ack_6060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2433_branch_ack_0, ack => timerDaemon_CP_5950_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_2432/do_while_stmt_2433/loop_taken/ack
      -- CP-element group 43: 	 branch_block_stmt_2432/do_while_stmt_2433/loop_taken/$exit
      -- 
    ack_6064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2433_branch_ack_1, ack => timerDaemon_CP_5950_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_2432/do_while_stmt_2433/$exit
      -- 
    timerDaemon_CP_5950_elements(44) <= timerDaemon_CP_5950_elements(3);
    timerDaemon_do_while_stmt_2433_terminator_6065: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_2433_terminator_6065", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_5950_elements(6),loop_continue => timerDaemon_CP_5950_elements(43),loop_terminate => timerDaemon_CP_5950_elements(42),loop_back => timerDaemon_CP_5950_elements(4),loop_exit => timerDaemon_CP_5950_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_2435_phi_seq_6023_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_5950_elements(21);
      timerDaemon_CP_5950_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_5950_elements(24);
      timerDaemon_CP_5950_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_5950_elements(26);
      timerDaemon_CP_5950_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_5950_elements(19);
      timerDaemon_CP_5950_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_5950_elements(30);
      timerDaemon_CP_5950_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_5950_elements(31);
      timerDaemon_CP_5950_elements(20) <= phi_mux_reqs(1);
      phi_stmt_2435_phi_seq_6023 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_2435_phi_seq_6023") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_5950_elements(11), 
          phi_sample_ack => timerDaemon_CP_5950_elements(17), 
          phi_update_req => timerDaemon_CP_5950_elements(13), 
          phi_update_ack => timerDaemon_CP_5950_elements(18), 
          phi_mux_ack => timerDaemon_CP_5950_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_5975_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_5950_elements(7);
        preds(1)  <= timerDaemon_CP_5950_elements(8);
        entry_tmerge_5975 : transition_merge -- 
          generic map(name => " entry_tmerge_5975")
          port map (preds => preds, symbol_out => timerDaemon_CP_5950_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_2435 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_2442_wire : std_logic_vector(0 downto 0);
    signal konst_2446_wire_constant : std_logic_vector(63 downto 0);
    signal konst_2454_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_2448 : std_logic_vector(63 downto 0);
    signal nCOUNTER_2448_2439_buffered : std_logic_vector(63 downto 0);
    signal req_2440 : std_logic_vector(0 downto 0);
    signal type_cast_2438_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_2446_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_2454_wire_constant <= "1";
    type_cast_2438_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_2435: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2438_wire_constant & nCOUNTER_2448_2439_buffered;
      req <= phi_stmt_2435_req_0 & phi_stmt_2435_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2435",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2435_ack_0,
          idata => idata,
          odata => COUNTER_2435,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2435
    nCOUNTER_2448_2439_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_2448_2439_buf_req_0;
      nCOUNTER_2448_2439_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_2448_2439_buf_req_1;
      nCOUNTER_2448_2439_buf_ack_1<= rack(0);
      nCOUNTER_2448_2439_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_2448_2439_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_2448,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_2448_2439_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_2440
    process(RPIPE_timer_req_2442_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_2442_wire(0 downto 0);
      req_2440 <= tmp_var; -- 
    end process;
    do_while_stmt_2433_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_2454_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2433_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2433_branch_req_0,
          ack0 => do_while_stmt_2433_branch_ack_0,
          ack1 => do_while_stmt_2433_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_2447_inst
    process(COUNTER_2435) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_2435, konst_2446_wire_constant, tmp_var);
      nCOUNTER_2448 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_2442_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_2442_inst_req_0;
      RPIPE_timer_req_2442_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_2442_inst_req_1;
      RPIPE_timer_req_2442_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_2442_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_2450_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_2450_inst_req_0;
      WPIPE_timer_resp_2450_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_2450_inst_req_1;
      WPIPE_timer_resp_2450_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_2440(0);
      data_in <= COUNTER_2435;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(2 downto 0);
  -- declarations related to module access_T
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      row_in : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      input_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module access_T
  signal access_T_row_in :  std_logic_vector(15 downto 0);
  signal access_T_chl_in :  std_logic_vector(15 downto 0);
  signal access_T_ct :  std_logic_vector(15 downto 0);
  signal access_T_in_args    : std_logic_vector(47 downto 0);
  signal access_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal access_T_tag_out   : std_logic_vector(1 downto 0);
  signal access_T_start_req : std_logic;
  signal access_T_start_ack : std_logic;
  signal access_T_fin_req   : std_logic;
  signal access_T_fin_ack : std_logic;
  -- caller side aggregated signals for module access_T
  signal access_T_call_reqs: std_logic_vector(0 downto 0);
  signal access_T_call_acks: std_logic_vector(0 downto 0);
  signal access_T_return_reqs: std_logic_vector(0 downto 0);
  signal access_T_return_acks: std_logic_vector(0 downto 0);
  signal access_T_call_data: std_logic_vector(47 downto 0);
  signal access_T_call_tag: std_logic_vector(0 downto 0);
  signal access_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module convolution3D
  component convolution3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      access_T_call_reqs : out  std_logic_vector(0 downto 0);
      access_T_call_acks : in   std_logic_vector(0 downto 0);
      access_T_call_data : out  std_logic_vector(47 downto 0);
      access_T_call_tag  :  out  std_logic_vector(0 downto 0);
      access_T_return_reqs : out  std_logic_vector(0 downto 0);
      access_T_return_acks : in   std_logic_vector(0 downto 0);
      access_T_return_tag :  in   std_logic_vector(0 downto 0);
      loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_call_data : out  std_logic_vector(79 downto 0);
      loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolution3D
  signal convolution3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolution3D_tag_out   : std_logic_vector(1 downto 0);
  signal convolution3D_start_req : std_logic;
  signal convolution3D_start_ack : std_logic;
  signal convolution3D_fin_req   : std_logic;
  signal convolution3D_fin_ack : std_logic;
  -- declarations related to module convolve
  component convolve is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe3_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      kernel_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_read_data : in   std_logic_vector(15 downto 0);
      kernel_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_read_data : in   std_logic_vector(15 downto 0);
      kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolve
  signal convolve_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolve_tag_out   : std_logic_vector(1 downto 0);
  signal convolve_start_req : std_logic;
  signal convolve_start_ack : std_logic;
  signal convolve_fin_req   : std_logic;
  signal convolve_fin_ack : std_logic;
  -- declarations related to module loadKernelChannel
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      num_chl : in  std_logic_vector(15 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_data : out  std_logic_vector(15 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadKernelChannel
  signal loadKernelChannel_start_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_num_chl :  std_logic_vector(15 downto 0);
  signal loadKernelChannel_in_args    : std_logic_vector(79 downto 0);
  signal loadKernelChannel_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadKernelChannel_tag_out   : std_logic_vector(1 downto 0);
  signal loadKernelChannel_start_req : std_logic;
  signal loadKernelChannel_start_ack : std_logic;
  signal loadKernelChannel_fin_req   : std_logic;
  signal loadKernelChannel_fin_ack : std_logic;
  -- caller side aggregated signals for module loadKernelChannel
  signal loadKernelChannel_call_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_data: std_logic_vector(79 downto 0);
  signal loadKernelChannel_call_tag: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe input_done_pipe
  signal input_done_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal input_done_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_done_pipe
  signal input_done_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_done_pipe_pipe_read_req: std_logic_vector(1 downto 0);
  signal input_done_pipe_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe input_pipe1
  signal input_pipe1_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe1
  signal input_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe2
  signal input_pipe2_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe2_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe2
  signal input_pipe2_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe2_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe3
  signal input_pipe3_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe3_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe3
  signal input_pipe3_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe3_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe1
  signal kernel_pipe1_pipe_write_data: std_logic_vector(15 downto 0);
  signal kernel_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe kernel_pipe1
  signal kernel_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe2
  signal kernel_pipe2_pipe_write_data: std_logic_vector(15 downto 0);
  signal kernel_pipe2_pipe_write_req: std_logic_vector(0 downto 0);
  signal kernel_pipe2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe kernel_pipe2
  signal kernel_pipe2_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe2_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe3
  signal kernel_pipe3_pipe_write_data: std_logic_vector(15 downto 0);
  signal kernel_pipe3_pipe_write_req: std_logic_vector(0 downto 0);
  signal kernel_pipe3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe kernel_pipe3
  signal kernel_pipe3_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe3_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe num_out_pipe
  signal num_out_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe num_out_pipe
  signal num_out_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe size_pipe
  signal size_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal size_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe size_pipe
  signal size_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal size_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module access_T
  access_T_row_in <= access_T_in_args(47 downto 32);
  access_T_chl_in <= access_T_in_args(31 downto 16);
  access_T_ct <= access_T_in_args(15 downto 0);
  -- call arbiter for module access_T
  access_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 48,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => access_T_call_reqs,
      call_acks => access_T_call_acks,
      return_reqs => access_T_return_reqs,
      return_acks => access_T_return_acks,
      call_data  => access_T_call_data,
      call_tag  => access_T_call_tag,
      return_tag  => access_T_return_tag,
      call_mtag => access_T_tag_in,
      return_mtag => access_T_tag_out,
      call_mreq => access_T_start_req,
      call_mack => access_T_start_ack,
      return_mreq => access_T_fin_req,
      return_mack => access_T_fin_ack,
      call_mdata => access_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  access_T_instance:access_T-- 
    generic map(tag_length => 2)
    port map(-- 
      row_in => access_T_row_in,
      chl_in => access_T_chl_in,
      ct => access_T_ct,
      start_req => access_T_start_req,
      start_ack => access_T_start_ack,
      fin_req => access_T_fin_req,
      fin_ack => access_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(19 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 0),
      input_pipe2_pipe_write_req => input_pipe2_pipe_write_req(0 downto 0),
      input_pipe2_pipe_write_ack => input_pipe2_pipe_write_ack(0 downto 0),
      input_pipe2_pipe_write_data => input_pipe2_pipe_write_data(15 downto 0),
      input_pipe3_pipe_write_req => input_pipe3_pipe_write_req(0 downto 0),
      input_pipe3_pipe_write_ack => input_pipe3_pipe_write_ack(0 downto 0),
      input_pipe3_pipe_write_data => input_pipe3_pipe_write_data(15 downto 0),
      input_pipe1_pipe_write_req => input_pipe1_pipe_write_req(0 downto 0),
      input_pipe1_pipe_write_ack => input_pipe1_pipe_write_ack(0 downto 0),
      input_pipe1_pipe_write_data => input_pipe1_pipe_write_data(15 downto 0),
      tag_in => access_T_tag_in,
      tag_out => access_T_tag_out-- 
    ); -- 
  -- module convolution3D
  convolution3D_instance:convolution3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolution3D_start_req,
      start_ack => convolution3D_start_ack,
      fin_req => convolution3D_fin_req,
      fin_ack => convolution3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(19 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(2 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(0 downto 0),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(0 downto 0),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(7 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(7 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(1 downto 1),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(1 downto 1),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(15 downto 8),
      num_out_pipe_pipe_write_req => num_out_pipe_pipe_write_req(0 downto 0),
      num_out_pipe_pipe_write_ack => num_out_pipe_pipe_write_ack(0 downto 0),
      num_out_pipe_pipe_write_data => num_out_pipe_pipe_write_data(15 downto 0),
      access_T_call_reqs => access_T_call_reqs(0 downto 0),
      access_T_call_acks => access_T_call_acks(0 downto 0),
      access_T_call_data => access_T_call_data(47 downto 0),
      access_T_call_tag => access_T_call_tag(0 downto 0),
      access_T_return_reqs => access_T_return_reqs(0 downto 0),
      access_T_return_acks => access_T_return_acks(0 downto 0),
      access_T_return_tag => access_T_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      loadKernelChannel_call_reqs => loadKernelChannel_call_reqs(0 downto 0),
      loadKernelChannel_call_acks => loadKernelChannel_call_acks(0 downto 0),
      loadKernelChannel_call_data => loadKernelChannel_call_data(79 downto 0),
      loadKernelChannel_call_tag => loadKernelChannel_call_tag(0 downto 0),
      loadKernelChannel_return_reqs => loadKernelChannel_return_reqs(0 downto 0),
      loadKernelChannel_return_acks => loadKernelChannel_return_acks(0 downto 0),
      loadKernelChannel_return_tag => loadKernelChannel_return_tag(0 downto 0),
      tag_in => convolution3D_tag_in,
      tag_out => convolution3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolution3D_tag_in <= (others => '0');
  convolution3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolution3D_start_req, start_ack => convolution3D_start_ack,  fin_req => convolution3D_fin_req,  fin_ack => convolution3D_fin_ack);
  -- module convolve
  convolve_instance:convolve-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolve_start_req,
      start_ack => convolve_start_ack,
      fin_req => convolve_fin_req,
      fin_ack => convolve_fin_ack,
      clk => clk,
      reset => reset,
      input_pipe2_pipe_read_req => input_pipe2_pipe_read_req(0 downto 0),
      input_pipe2_pipe_read_ack => input_pipe2_pipe_read_ack(0 downto 0),
      input_pipe2_pipe_read_data => input_pipe2_pipe_read_data(15 downto 0),
      input_pipe3_pipe_read_req => input_pipe3_pipe_read_req(0 downto 0),
      input_pipe3_pipe_read_ack => input_pipe3_pipe_read_ack(0 downto 0),
      input_pipe3_pipe_read_data => input_pipe3_pipe_read_data(15 downto 0),
      input_pipe1_pipe_read_req => input_pipe1_pipe_read_req(0 downto 0),
      input_pipe1_pipe_read_ack => input_pipe1_pipe_read_ack(0 downto 0),
      input_pipe1_pipe_read_data => input_pipe1_pipe_read_data(15 downto 0),
      kernel_pipe2_pipe_read_req => kernel_pipe2_pipe_read_req(0 downto 0),
      kernel_pipe2_pipe_read_ack => kernel_pipe2_pipe_read_ack(0 downto 0),
      kernel_pipe2_pipe_read_data => kernel_pipe2_pipe_read_data(15 downto 0),
      kernel_pipe3_pipe_read_req => kernel_pipe3_pipe_read_req(0 downto 0),
      kernel_pipe3_pipe_read_ack => kernel_pipe3_pipe_read_ack(0 downto 0),
      kernel_pipe3_pipe_read_data => kernel_pipe3_pipe_read_data(15 downto 0),
      kernel_pipe1_pipe_read_req => kernel_pipe1_pipe_read_req(0 downto 0),
      kernel_pipe1_pipe_read_ack => kernel_pipe1_pipe_read_ack(0 downto 0),
      kernel_pipe1_pipe_read_data => kernel_pipe1_pipe_read_data(15 downto 0),
      num_out_pipe_pipe_read_req => num_out_pipe_pipe_read_req(0 downto 0),
      num_out_pipe_pipe_read_ack => num_out_pipe_pipe_read_ack(0 downto 0),
      num_out_pipe_pipe_read_data => num_out_pipe_pipe_read_data(15 downto 0),
      size_pipe_pipe_read_req => size_pipe_pipe_read_req(0 downto 0),
      size_pipe_pipe_read_ack => size_pipe_pipe_read_ack(0 downto 0),
      size_pipe_pipe_read_data => size_pipe_pipe_read_data(15 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(0 downto 0),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(0 downto 0),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(7 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(7 downto 0),
      tag_in => convolve_tag_in,
      tag_out => convolve_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolve_tag_in <= (others => '0');
  convolve_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolve_start_req, start_ack => convolve_start_ack,  fin_req => convolve_fin_req,  fin_ack => convolve_fin_ack);
  -- module loadKernelChannel
  loadKernelChannel_start_add <= loadKernelChannel_in_args(79 downto 16);
  loadKernelChannel_num_chl <= loadKernelChannel_in_args(15 downto 0);
  -- call arbiter for module loadKernelChannel
  loadKernelChannel_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 80,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadKernelChannel_call_reqs,
      call_acks => loadKernelChannel_call_acks,
      return_reqs => loadKernelChannel_return_reqs,
      return_acks => loadKernelChannel_return_acks,
      call_data  => loadKernelChannel_call_data,
      call_tag  => loadKernelChannel_call_tag,
      return_tag  => loadKernelChannel_return_tag,
      call_mtag => loadKernelChannel_tag_in,
      return_mtag => loadKernelChannel_tag_out,
      call_mreq => loadKernelChannel_start_req,
      call_mack => loadKernelChannel_start_ack,
      return_mreq => loadKernelChannel_fin_req,
      return_mack => loadKernelChannel_fin_ack,
      call_mdata => loadKernelChannel_in_args,
      clk => clk, 
      reset => reset --
    ); --
  loadKernelChannel_instance:loadKernelChannel-- 
    generic map(tag_length => 2)
    port map(-- 
      start_add => loadKernelChannel_start_add,
      num_chl => loadKernelChannel_num_chl,
      start_req => loadKernelChannel_start_req,
      start_ack => loadKernelChannel_start_ack,
      fin_req => loadKernelChannel_fin_req,
      fin_ack => loadKernelChannel_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(1 downto 1),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(1 downto 1),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(15 downto 8),
      kernel_pipe2_pipe_write_req => kernel_pipe2_pipe_write_req(0 downto 0),
      kernel_pipe2_pipe_write_ack => kernel_pipe2_pipe_write_ack(0 downto 0),
      kernel_pipe2_pipe_write_data => kernel_pipe2_pipe_write_data(15 downto 0),
      kernel_pipe3_pipe_write_req => kernel_pipe3_pipe_write_req(0 downto 0),
      kernel_pipe3_pipe_write_ack => kernel_pipe3_pipe_write_ack(0 downto 0),
      kernel_pipe3_pipe_write_data => kernel_pipe3_pipe_write_data(15 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(0 downto 0),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(0 downto 0),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(15 downto 0),
      size_pipe_pipe_write_req => size_pipe_pipe_write_req(0 downto 0),
      size_pipe_pipe_write_ack => size_pipe_pipe_write_ack(0 downto 0),
      size_pipe_pipe_write_data => size_pipe_pipe_write_data(15 downto 0),
      tag_in => loadKernelChannel_tag_in,
      tag_out => loadKernelChannel_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  input_done_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_done_pipe",
      num_reads => 2,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => input_done_pipe_pipe_read_req,
      read_ack => input_done_pipe_pipe_read_ack,
      read_data => input_done_pipe_pipe_read_data,
      write_req => input_done_pipe_pipe_write_req,
      write_ack => input_done_pipe_pipe_write_ack,
      write_data => input_done_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe1_pipe_read_req,
      read_ack => input_pipe1_pipe_read_ack,
      read_data => input_pipe1_pipe_read_data,
      write_req => input_pipe1_pipe_write_req,
      write_ack => input_pipe1_pipe_write_ack,
      write_data => input_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe2",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe2_pipe_read_req,
      read_ack => input_pipe2_pipe_read_ack,
      read_data => input_pipe2_pipe_read_data,
      write_req => input_pipe2_pipe_write_req,
      write_ack => input_pipe2_pipe_write_ack,
      write_data => input_pipe2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe3",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => input_pipe3_pipe_read_req,
      read_ack => input_pipe3_pipe_read_ack,
      read_data => input_pipe3_pipe_read_data,
      write_req => input_pipe3_pipe_write_req,
      write_ack => input_pipe3_pipe_write_ack,
      write_data => input_pipe3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => kernel_pipe1_pipe_read_req,
      read_ack => kernel_pipe1_pipe_read_ack,
      read_data => kernel_pipe1_pipe_read_data,
      write_req => kernel_pipe1_pipe_write_req,
      write_ack => kernel_pipe1_pipe_write_ack,
      write_data => kernel_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe2",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => kernel_pipe2_pipe_read_req,
      read_ack => kernel_pipe2_pipe_read_ack,
      read_data => kernel_pipe2_pipe_read_data,
      write_req => kernel_pipe2_pipe_write_req,
      write_ack => kernel_pipe2_pipe_write_ack,
      write_data => kernel_pipe2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe3",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 400 --
    )
    port map( -- 
      read_req => kernel_pipe3_pipe_read_req,
      read_ack => kernel_pipe3_pipe_read_ack,
      read_data => kernel_pipe3_pipe_read_data,
      write_req => kernel_pipe3_pipe_write_req,
      write_ack => kernel_pipe3_pipe_write_ack,
      write_data => kernel_pipe3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  num_out_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe num_out_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => num_out_pipe_pipe_read_req,
      read_ack => num_out_pipe_pipe_read_ack,
      read_data => num_out_pipe_pipe_read_data,
      write_req => num_out_pipe_pipe_write_req,
      write_ack => num_out_pipe_pipe_write_ack,
      write_data => num_out_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  size_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe size_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 11 --
    )
    port map( -- 
      read_req => size_pipe_pipe_read_req,
      read_ack => size_pipe_pipe_read_ack,
      read_data => size_pipe_pipe_read_data,
      write_req => size_pipe_pipe_write_req,
      write_ack => size_pipe_pipe_write_ack,
      write_data => size_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
