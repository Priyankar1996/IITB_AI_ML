-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(31 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(31 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(31 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(31 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(31 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(31 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(31 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(31 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_39_start: Boolean;
  signal convTranspose_CP_39_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_735_inst_req_0 : boolean;
  signal type_cast_528_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1002_inst_ack_1 : boolean;
  signal type_cast_735_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_749_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1002_inst_req_0 : boolean;
  signal type_cast_528_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1062_inst_ack_1 : boolean;
  signal type_cast_735_inst_req_1 : boolean;
  signal if_stmt_604_branch_ack_1 : boolean;
  signal type_cast_717_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_749_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_542_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_542_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1023_inst_ack_1 : boolean;
  signal type_cast_474_inst_req_1 : boolean;
  signal type_cast_717_inst_req_1 : boolean;
  signal ptr_deref_590_store_0_req_1 : boolean;
  signal type_cast_1162_inst_req_0 : boolean;
  signal type_cast_735_inst_ack_0 : boolean;
  signal type_cast_717_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_749_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_749_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1071_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1011_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_488_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_488_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_488_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_488_inst_req_0 : boolean;
  signal type_cast_528_inst_ack_1 : boolean;
  signal type_cast_528_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_993_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 : boolean;
  signal type_cast_717_inst_req_0 : boolean;
  signal WPIPE_Block1_start_993_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_560_inst_ack_1 : boolean;
  signal type_cast_38_inst_req_0 : boolean;
  signal type_cast_38_inst_ack_0 : boolean;
  signal type_cast_38_inst_req_1 : boolean;
  signal type_cast_38_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_664_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_134_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_47_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_560_inst_req_1 : boolean;
  signal type_cast_51_inst_req_0 : boolean;
  signal type_cast_51_inst_ack_0 : boolean;
  signal type_cast_51_inst_req_1 : boolean;
  signal type_cast_51_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1038_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_59_inst_ack_1 : boolean;
  signal type_cast_681_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_524_inst_ack_0 : boolean;
  signal type_cast_63_inst_req_0 : boolean;
  signal type_cast_63_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1005_inst_ack_0 : boolean;
  signal type_cast_63_inst_req_1 : boolean;
  signal type_cast_63_inst_ack_1 : boolean;
  signal if_stmt_604_branch_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_524_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_72_inst_ack_1 : boolean;
  signal type_cast_681_inst_req_1 : boolean;
  signal ptr_deref_590_store_0_ack_0 : boolean;
  signal type_cast_76_inst_req_0 : boolean;
  signal type_cast_76_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1038_inst_req_1 : boolean;
  signal type_cast_76_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1011_inst_req_1 : boolean;
  signal type_cast_76_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_524_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_req_0 : boolean;
  signal type_cast_582_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_664_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_84_inst_ack_1 : boolean;
  signal type_cast_681_inst_ack_0 : boolean;
  signal type_cast_681_inst_req_0 : boolean;
  signal array_obj_ref_660_index_offset_ack_1 : boolean;
  signal WPIPE_Block2_start_1029_inst_req_0 : boolean;
  signal ptr_deref_590_store_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_560_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1005_inst_req_0 : boolean;
  signal type_cast_88_inst_req_0 : boolean;
  signal type_cast_582_inst_req_1 : boolean;
  signal type_cast_88_inst_ack_0 : boolean;
  signal type_cast_88_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1050_inst_req_0 : boolean;
  signal type_cast_88_inst_ack_1 : boolean;
  signal type_cast_1162_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_97_inst_ack_1 : boolean;
  signal array_obj_ref_660_index_offset_req_1 : boolean;
  signal WPIPE_Block1_start_987_inst_req_1 : boolean;
  signal type_cast_101_inst_req_0 : boolean;
  signal type_cast_101_inst_ack_0 : boolean;
  signal type_cast_101_inst_req_1 : boolean;
  signal type_cast_101_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_524_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_664_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_req_0 : boolean;
  signal type_cast_582_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_109_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1071_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_560_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1029_inst_ack_0 : boolean;
  signal type_cast_113_inst_req_0 : boolean;
  signal type_cast_582_inst_req_0 : boolean;
  signal type_cast_113_inst_ack_0 : boolean;
  signal type_cast_113_inst_req_1 : boolean;
  signal type_cast_113_inst_ack_1 : boolean;
  signal type_cast_699_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_122_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_987_inst_ack_1 : boolean;
  signal array_obj_ref_660_index_offset_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_695_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1005_inst_req_1 : boolean;
  signal array_obj_ref_660_index_offset_req_0 : boolean;
  signal type_cast_126_inst_req_0 : boolean;
  signal type_cast_126_inst_ack_0 : boolean;
  signal type_cast_126_inst_req_1 : boolean;
  signal type_cast_126_inst_ack_1 : boolean;
  signal type_cast_699_inst_req_1 : boolean;
  signal WPIPE_Block1_start_990_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1026_inst_req_0 : boolean;
  signal type_cast_361_inst_req_0 : boolean;
  signal type_cast_361_inst_ack_0 : boolean;
  signal type_cast_361_inst_req_1 : boolean;
  signal type_cast_361_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1059_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_370_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_370_inst_ack_0 : boolean;
  signal type_cast_492_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_370_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_370_inst_ack_1 : boolean;
  signal type_cast_138_inst_req_0 : boolean;
  signal type_cast_138_inst_ack_0 : boolean;
  signal type_cast_138_inst_req_1 : boolean;
  signal type_cast_138_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_731_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1011_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_ack_0 : boolean;
  signal type_cast_510_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_664_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_147_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_695_inst_req_1 : boolean;
  signal type_cast_151_inst_req_0 : boolean;
  signal type_cast_151_inst_ack_0 : boolean;
  signal type_cast_151_inst_req_1 : boolean;
  signal WPIPE_Block1_start_996_inst_req_0 : boolean;
  signal type_cast_151_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1068_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_731_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1074_inst_req_1 : boolean;
  signal type_cast_510_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1050_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_159_inst_ack_1 : boolean;
  signal type_cast_492_inst_ack_1 : boolean;
  signal type_cast_163_inst_req_0 : boolean;
  signal type_cast_163_inst_ack_0 : boolean;
  signal type_cast_163_inst_req_1 : boolean;
  signal type_cast_163_inst_ack_1 : boolean;
  signal type_cast_699_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_172_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_677_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1026_inst_req_1 : boolean;
  signal type_cast_176_inst_req_0 : boolean;
  signal type_cast_176_inst_ack_0 : boolean;
  signal type_cast_176_inst_req_1 : boolean;
  signal type_cast_176_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1074_inst_ack_1 : boolean;
  signal addr_of_661_final_reg_ack_1 : boolean;
  signal type_cast_510_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1005_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_ack_0 : boolean;
  signal type_cast_510_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_184_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_713_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_677_inst_req_1 : boolean;
  signal type_cast_188_inst_req_0 : boolean;
  signal type_cast_188_inst_ack_0 : boolean;
  signal type_cast_188_inst_req_1 : boolean;
  signal type_cast_188_inst_ack_1 : boolean;
  signal type_cast_699_inst_req_0 : boolean;
  signal addr_of_661_final_reg_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_731_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_578_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_197_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_713_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_677_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_695_inst_ack_0 : boolean;
  signal type_cast_201_inst_req_0 : boolean;
  signal type_cast_201_inst_ack_0 : boolean;
  signal type_cast_201_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_578_inst_req_1 : boolean;
  signal type_cast_201_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_731_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_257_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_257_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_257_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_257_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_677_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1029_inst_req_1 : boolean;
  signal type_cast_631_inst_ack_1 : boolean;
  signal type_cast_261_inst_req_0 : boolean;
  signal type_cast_261_inst_ack_0 : boolean;
  signal type_cast_261_inst_req_1 : boolean;
  signal type_cast_261_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1029_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1002_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_270_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_578_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_270_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_270_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_270_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_695_inst_req_0 : boolean;
  signal type_cast_631_inst_req_1 : boolean;
  signal type_cast_274_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_578_inst_req_0 : boolean;
  signal type_cast_274_inst_ack_0 : boolean;
  signal type_cast_274_inst_req_1 : boolean;
  signal type_cast_274_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_506_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_282_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_282_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_506_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_282_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_282_inst_ack_1 : boolean;
  signal type_cast_286_inst_req_0 : boolean;
  signal type_cast_286_inst_ack_0 : boolean;
  signal type_cast_286_inst_req_1 : boolean;
  signal type_cast_286_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_990_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_295_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_295_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_295_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_295_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_713_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1071_inst_ack_1 : boolean;
  signal type_cast_546_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1026_inst_ack_0 : boolean;
  signal type_cast_299_inst_req_0 : boolean;
  signal type_cast_299_inst_ack_0 : boolean;
  signal type_cast_631_inst_ack_0 : boolean;
  signal type_cast_299_inst_req_1 : boolean;
  signal type_cast_299_inst_ack_1 : boolean;
  signal addr_of_661_final_reg_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_506_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_307_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_307_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_506_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_307_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_307_inst_ack_1 : boolean;
  signal type_cast_546_inst_req_1 : boolean;
  signal type_cast_311_inst_req_0 : boolean;
  signal type_cast_311_inst_ack_0 : boolean;
  signal type_cast_631_inst_req_0 : boolean;
  signal type_cast_311_inst_req_1 : boolean;
  signal type_cast_311_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_320_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1050_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_320_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_320_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_320_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_713_inst_req_0 : boolean;
  signal type_cast_668_inst_ack_1 : boolean;
  signal type_cast_324_inst_req_0 : boolean;
  signal type_cast_324_inst_ack_0 : boolean;
  signal type_cast_324_inst_req_1 : boolean;
  signal type_cast_324_inst_ack_1 : boolean;
  signal addr_of_661_final_reg_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_332_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_332_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_332_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_332_inst_ack_1 : boolean;
  signal type_cast_668_inst_req_1 : boolean;
  signal type_cast_336_inst_req_0 : boolean;
  signal type_cast_336_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1038_inst_ack_1 : boolean;
  signal type_cast_336_inst_req_1 : boolean;
  signal type_cast_336_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1002_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_345_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_345_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_990_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_345_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_345_inst_ack_1 : boolean;
  signal type_cast_668_inst_ack_0 : boolean;
  signal type_cast_546_inst_ack_0 : boolean;
  signal type_cast_349_inst_req_0 : boolean;
  signal type_cast_349_inst_ack_0 : boolean;
  signal type_cast_349_inst_req_1 : boolean;
  signal type_cast_564_inst_ack_1 : boolean;
  signal type_cast_349_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1077_inst_req_0 : boolean;
  signal type_cast_492_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_357_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1050_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_357_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_357_inst_req_1 : boolean;
  signal type_cast_564_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_357_inst_ack_1 : boolean;
  signal type_cast_668_inst_req_0 : boolean;
  signal type_cast_546_inst_req_0 : boolean;
  signal type_cast_374_inst_req_0 : boolean;
  signal type_cast_564_inst_ack_0 : boolean;
  signal type_cast_374_inst_ack_0 : boolean;
  signal type_cast_374_inst_req_1 : boolean;
  signal type_cast_374_inst_ack_1 : boolean;
  signal type_cast_492_inst_req_0 : boolean;
  signal if_stmt_604_branch_ack_0 : boolean;
  signal ptr_deref_590_store_0_ack_1 : boolean;
  signal WPIPE_Block2_start_1026_inst_ack_1 : boolean;
  signal if_stmt_388_branch_req_0 : boolean;
  signal if_stmt_388_branch_ack_1 : boolean;
  signal type_cast_474_inst_ack_1 : boolean;
  signal if_stmt_388_branch_ack_0 : boolean;
  signal type_cast_564_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1041_inst_req_0 : boolean;
  signal if_stmt_403_branch_req_0 : boolean;
  signal WPIPE_Block2_start_1032_inst_req_1 : boolean;
  signal WPIPE_Block1_start_996_inst_ack_0 : boolean;
  signal if_stmt_403_branch_ack_1 : boolean;
  signal if_stmt_403_branch_ack_0 : boolean;
  signal WPIPE_Block2_start_1041_inst_ack_0 : boolean;
  signal type_cast_424_inst_req_0 : boolean;
  signal type_cast_424_inst_ack_0 : boolean;
  signal type_cast_424_inst_req_1 : boolean;
  signal type_cast_424_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_542_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_542_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1011_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1032_inst_req_0 : boolean;
  signal array_obj_ref_453_index_offset_req_0 : boolean;
  signal WPIPE_Block2_start_1032_inst_ack_0 : boolean;
  signal array_obj_ref_453_index_offset_ack_0 : boolean;
  signal array_obj_ref_453_index_offset_req_1 : boolean;
  signal array_obj_ref_453_index_offset_ack_1 : boolean;
  signal addr_of_454_final_reg_req_0 : boolean;
  signal addr_of_454_final_reg_ack_0 : boolean;
  signal addr_of_454_final_reg_req_1 : boolean;
  signal addr_of_454_final_reg_ack_1 : boolean;
  signal WPIPE_Block3_start_1059_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_457_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_457_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1008_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_457_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_457_inst_ack_1 : boolean;
  signal type_cast_461_inst_req_0 : boolean;
  signal type_cast_461_inst_ack_0 : boolean;
  signal type_cast_461_inst_req_1 : boolean;
  signal type_cast_461_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_470_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_470_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_470_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_470_inst_ack_1 : boolean;
  signal type_cast_474_inst_req_0 : boolean;
  signal type_cast_474_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1023_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1062_inst_req_1 : boolean;
  signal type_cast_753_inst_req_0 : boolean;
  signal type_cast_753_inst_ack_0 : boolean;
  signal type_cast_753_inst_req_1 : boolean;
  signal type_cast_753_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_767_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_767_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_767_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_767_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1071_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1065_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1053_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1023_inst_ack_0 : boolean;
  signal type_cast_771_inst_req_0 : boolean;
  signal type_cast_771_inst_ack_0 : boolean;
  signal type_cast_771_inst_req_1 : boolean;
  signal type_cast_1162_inst_req_1 : boolean;
  signal type_cast_771_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1068_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1053_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1056_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1056_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_785_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1047_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_785_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_785_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_785_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1023_inst_req_0 : boolean;
  signal type_cast_789_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1047_inst_req_1 : boolean;
  signal type_cast_789_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1062_inst_ack_0 : boolean;
  signal type_cast_789_inst_req_1 : boolean;
  signal type_cast_1162_inst_ack_1 : boolean;
  signal type_cast_789_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1074_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1077_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1068_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1053_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1053_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1068_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1038_inst_req_0 : boolean;
  signal ptr_deref_797_store_0_req_0 : boolean;
  signal ptr_deref_797_store_0_ack_0 : boolean;
  signal ptr_deref_797_store_0_req_1 : boolean;
  signal ptr_deref_797_store_0_ack_1 : boolean;
  signal WPIPE_Block3_start_1077_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1059_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1020_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1062_inst_req_0 : boolean;
  signal WPIPE_Block1_start_993_inst_ack_0 : boolean;
  signal if_stmt_811_branch_req_0 : boolean;
  signal WPIPE_Block3_start_1065_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1020_inst_req_1 : boolean;
  signal WPIPE_Block1_start_993_inst_req_0 : boolean;
  signal if_stmt_811_branch_ack_1 : boolean;
  signal if_stmt_811_branch_ack_0 : boolean;
  signal WPIPE_Block2_start_1008_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1074_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1035_inst_ack_1 : boolean;
  signal if_stmt_836_branch_req_0 : boolean;
  signal WPIPE_Block2_start_1035_inst_req_1 : boolean;
  signal if_stmt_836_branch_ack_1 : boolean;
  signal if_stmt_836_branch_ack_0 : boolean;
  signal WPIPE_Block3_start_1056_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1008_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1035_inst_ack_0 : boolean;
  signal type_cast_863_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1047_inst_ack_0 : boolean;
  signal type_cast_863_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1035_inst_req_0 : boolean;
  signal type_cast_863_inst_req_1 : boolean;
  signal type_cast_863_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1059_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1020_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_990_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1020_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1056_inst_req_0 : boolean;
  signal array_obj_ref_892_index_offset_req_0 : boolean;
  signal WPIPE_Block3_start_1047_inst_req_0 : boolean;
  signal array_obj_ref_892_index_offset_ack_0 : boolean;
  signal array_obj_ref_892_index_offset_req_1 : boolean;
  signal array_obj_ref_892_index_offset_ack_1 : boolean;
  signal addr_of_893_final_reg_req_0 : boolean;
  signal addr_of_893_final_reg_ack_0 : boolean;
  signal addr_of_893_final_reg_req_1 : boolean;
  signal addr_of_893_final_reg_ack_1 : boolean;
  signal WPIPE_Block1_start_999_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1017_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1017_inst_req_1 : boolean;
  signal WPIPE_Block1_start_999_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1017_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1017_inst_req_0 : boolean;
  signal WPIPE_Block1_start_987_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1044_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1044_inst_req_1 : boolean;
  signal ptr_deref_896_store_0_req_0 : boolean;
  signal ptr_deref_896_store_0_ack_0 : boolean;
  signal WPIPE_Block1_start_987_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1008_inst_ack_0 : boolean;
  signal ptr_deref_896_store_0_req_1 : boolean;
  signal ptr_deref_896_store_0_ack_1 : boolean;
  signal WPIPE_Block1_start_999_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_999_inst_req_0 : boolean;
  signal if_stmt_911_branch_req_0 : boolean;
  signal WPIPE_Block2_start_1014_inst_ack_1 : boolean;
  signal if_stmt_911_branch_ack_1 : boolean;
  signal if_stmt_911_branch_ack_0 : boolean;
  signal WPIPE_Block2_start_1014_inst_req_1 : boolean;
  signal call_stmt_922_call_req_0 : boolean;
  signal WPIPE_Block2_start_1044_inst_ack_0 : boolean;
  signal call_stmt_922_call_ack_0 : boolean;
  signal WPIPE_Block2_start_1032_inst_ack_1 : boolean;
  signal if_stmt_1287_branch_ack_1 : boolean;
  signal call_stmt_922_call_req_1 : boolean;
  signal WPIPE_Block2_start_1044_inst_req_0 : boolean;
  signal call_stmt_922_call_ack_1 : boolean;
  signal type_cast_927_inst_req_0 : boolean;
  signal type_cast_927_inst_ack_0 : boolean;
  signal type_cast_927_inst_req_1 : boolean;
  signal type_cast_927_inst_ack_1 : boolean;
  signal if_stmt_1287_branch_ack_0 : boolean;
  signal WPIPE_Block2_start_1014_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_929_inst_req_0 : boolean;
  signal WPIPE_Block0_start_929_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_929_inst_req_1 : boolean;
  signal WPIPE_Block0_start_929_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1065_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1065_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1014_inst_req_0 : boolean;
  signal WPIPE_Block0_start_932_inst_req_0 : boolean;
  signal WPIPE_Block0_start_932_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_932_inst_req_1 : boolean;
  signal WPIPE_Block2_start_1041_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_932_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_996_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_935_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1041_inst_req_1 : boolean;
  signal WPIPE_Block0_start_935_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_996_inst_req_1 : boolean;
  signal WPIPE_Block0_start_935_inst_req_1 : boolean;
  signal WPIPE_Block0_start_935_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_938_inst_req_0 : boolean;
  signal WPIPE_Block0_start_938_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_938_inst_req_1 : boolean;
  signal WPIPE_Block0_start_938_inst_ack_1 : boolean;
  signal type_cast_447_inst_req_0 : boolean;
  signal phi_stmt_1159_req_0 : boolean;
  signal WPIPE_Block0_start_941_inst_req_0 : boolean;
  signal WPIPE_Block0_start_941_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_941_inst_req_1 : boolean;
  signal WPIPE_Block0_start_941_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_944_inst_req_0 : boolean;
  signal WPIPE_Block0_start_944_inst_ack_0 : boolean;
  signal type_cast_447_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_944_inst_req_1 : boolean;
  signal WPIPE_Block0_start_944_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_947_inst_req_0 : boolean;
  signal WPIPE_Block0_start_947_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_947_inst_req_1 : boolean;
  signal WPIPE_Block0_start_947_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_950_inst_req_0 : boolean;
  signal phi_stmt_1159_ack_0 : boolean;
  signal WPIPE_Block0_start_950_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_950_inst_req_1 : boolean;
  signal WPIPE_Block0_start_950_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_953_inst_req_0 : boolean;
  signal WPIPE_Block0_start_953_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1077_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_953_inst_req_1 : boolean;
  signal WPIPE_Block0_start_953_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_956_inst_req_0 : boolean;
  signal WPIPE_Block0_start_956_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_956_inst_req_1 : boolean;
  signal WPIPE_Block0_start_956_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_960_inst_req_0 : boolean;
  signal WPIPE_Block0_start_960_inst_ack_0 : boolean;
  signal type_cast_447_inst_req_1 : boolean;
  signal WPIPE_Block0_start_960_inst_req_1 : boolean;
  signal WPIPE_Block0_start_960_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_963_inst_req_0 : boolean;
  signal WPIPE_Block0_start_963_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_963_inst_req_1 : boolean;
  signal WPIPE_Block0_start_963_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_966_inst_req_0 : boolean;
  signal WPIPE_Block0_start_966_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_966_inst_req_1 : boolean;
  signal WPIPE_Block0_start_966_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_969_inst_req_0 : boolean;
  signal WPIPE_Block1_start_969_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_969_inst_req_1 : boolean;
  signal WPIPE_Block1_start_969_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_972_inst_req_0 : boolean;
  signal WPIPE_Block1_start_972_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_972_inst_req_1 : boolean;
  signal WPIPE_Block1_start_972_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_975_inst_req_0 : boolean;
  signal WPIPE_Block1_start_975_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_975_inst_req_1 : boolean;
  signal WPIPE_Block1_start_975_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_978_inst_req_0 : boolean;
  signal WPIPE_Block1_start_978_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_978_inst_req_1 : boolean;
  signal WPIPE_Block1_start_978_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_981_inst_req_0 : boolean;
  signal WPIPE_Block1_start_981_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_981_inst_req_1 : boolean;
  signal WPIPE_Block1_start_981_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_984_inst_req_0 : boolean;
  signal WPIPE_Block1_start_984_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_984_inst_req_1 : boolean;
  signal WPIPE_Block1_start_984_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1080_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1080_inst_ack_0 : boolean;
  signal phi_stmt_441_req_0 : boolean;
  signal WPIPE_Block3_start_1080_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1080_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1083_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1083_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1083_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1083_inst_ack_1 : boolean;
  signal RPIPE_Block0_done_1087_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1087_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1087_inst_req_1 : boolean;
  signal phi_stmt_1159_req_1 : boolean;
  signal RPIPE_Block0_done_1087_inst_ack_1 : boolean;
  signal phi_stmt_648_ack_0 : boolean;
  signal RPIPE_Block1_done_1090_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1090_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1090_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1090_inst_ack_1 : boolean;
  signal RPIPE_Block2_done_1093_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1093_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1093_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1093_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1096_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1096_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1096_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1096_inst_ack_1 : boolean;
  signal phi_stmt_648_req_0 : boolean;
  signal call_stmt_1100_call_req_0 : boolean;
  signal call_stmt_1100_call_ack_0 : boolean;
  signal call_stmt_1100_call_req_1 : boolean;
  signal call_stmt_1100_call_ack_1 : boolean;
  signal type_cast_651_inst_ack_1 : boolean;
  signal if_stmt_1287_branch_req_0 : boolean;
  signal type_cast_1104_inst_req_0 : boolean;
  signal type_cast_1104_inst_ack_0 : boolean;
  signal type_cast_1104_inst_req_1 : boolean;
  signal type_cast_1104_inst_ack_1 : boolean;
  signal type_cast_651_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1111_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1111_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1111_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1111_inst_ack_1 : boolean;
  signal type_cast_651_inst_ack_0 : boolean;
  signal type_cast_651_inst_req_0 : boolean;
  signal if_stmt_1115_branch_req_0 : boolean;
  signal if_stmt_1115_branch_ack_1 : boolean;
  signal if_stmt_1115_branch_ack_0 : boolean;
  signal phi_stmt_441_ack_0 : boolean;
  signal type_cast_1142_inst_req_0 : boolean;
  signal type_cast_1142_inst_ack_0 : boolean;
  signal type_cast_1142_inst_req_1 : boolean;
  signal type_cast_1142_inst_ack_1 : boolean;
  signal array_obj_ref_1171_index_offset_req_0 : boolean;
  signal array_obj_ref_1171_index_offset_ack_0 : boolean;
  signal array_obj_ref_1171_index_offset_req_1 : boolean;
  signal array_obj_ref_1171_index_offset_ack_1 : boolean;
  signal addr_of_1172_final_reg_req_0 : boolean;
  signal addr_of_1172_final_reg_ack_0 : boolean;
  signal addr_of_1172_final_reg_req_1 : boolean;
  signal addr_of_1172_final_reg_ack_1 : boolean;
  signal phi_stmt_441_req_1 : boolean;
  signal ptr_deref_1176_load_0_req_0 : boolean;
  signal ptr_deref_1176_load_0_ack_0 : boolean;
  signal phi_stmt_880_req_1 : boolean;
  signal type_cast_447_inst_ack_1 : boolean;
  signal ptr_deref_1176_load_0_req_1 : boolean;
  signal phi_stmt_648_req_1 : boolean;
  signal ptr_deref_1176_load_0_ack_1 : boolean;
  signal type_cast_1180_inst_req_0 : boolean;
  signal type_cast_1180_inst_ack_0 : boolean;
  signal type_cast_1180_inst_req_1 : boolean;
  signal type_cast_1180_inst_ack_1 : boolean;
  signal type_cast_1190_inst_req_0 : boolean;
  signal type_cast_1190_inst_ack_0 : boolean;
  signal type_cast_1190_inst_req_1 : boolean;
  signal type_cast_1190_inst_ack_1 : boolean;
  signal type_cast_1200_inst_req_0 : boolean;
  signal type_cast_1200_inst_ack_0 : boolean;
  signal type_cast_1200_inst_req_1 : boolean;
  signal phi_stmt_880_ack_0 : boolean;
  signal type_cast_1200_inst_ack_1 : boolean;
  signal type_cast_1210_inst_req_0 : boolean;
  signal type_cast_1210_inst_ack_0 : boolean;
  signal type_cast_1210_inst_req_1 : boolean;
  signal phi_stmt_880_req_0 : boolean;
  signal type_cast_1210_inst_ack_1 : boolean;
  signal type_cast_883_inst_ack_1 : boolean;
  signal type_cast_1220_inst_req_0 : boolean;
  signal type_cast_883_inst_req_1 : boolean;
  signal type_cast_1220_inst_ack_0 : boolean;
  signal type_cast_1220_inst_req_1 : boolean;
  signal type_cast_1220_inst_ack_1 : boolean;
  signal type_cast_1230_inst_req_0 : boolean;
  signal type_cast_883_inst_ack_0 : boolean;
  signal type_cast_1230_inst_ack_0 : boolean;
  signal type_cast_1230_inst_req_1 : boolean;
  signal type_cast_883_inst_req_0 : boolean;
  signal type_cast_1230_inst_ack_1 : boolean;
  signal type_cast_1240_inst_req_0 : boolean;
  signal type_cast_1240_inst_ack_0 : boolean;
  signal type_cast_1240_inst_req_1 : boolean;
  signal type_cast_1240_inst_ack_1 : boolean;
  signal type_cast_1250_inst_req_0 : boolean;
  signal type_cast_1250_inst_ack_0 : boolean;
  signal type_cast_1250_inst_req_1 : boolean;
  signal type_cast_1250_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1252_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1252_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1252_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1252_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1255_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1255_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1255_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1255_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1258_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1258_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1258_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1258_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1261_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1261_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1261_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1261_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1264_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1264_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1264_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1264_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1267_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1267_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1267_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1267_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1270_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1270_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1270_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1270_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1273_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1273_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1273_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1273_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_39_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_39_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_39: Block -- control-path 
    signal convTranspose_CP_39_elements: BooleanArray(405 downto 0);
    -- 
  begin -- 
    convTranspose_CP_39_elements(0) <= convTranspose_CP_39_start;
    convTranspose_CP_39_symbol <= convTranspose_CP_39_elements(405);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	84 
    -- CP-element group 0: 	88 
    -- CP-element group 0: 	80 
    -- CP-element group 0: 	92 
    -- CP-element group 0: 	96 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	72 
    -- CP-element group 0: 	76 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	64 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0:  members (80) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_32/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/branch_block_stmt_32__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_34_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_34_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_34_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_38_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_38_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_38_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_138_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_51_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_51_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_51_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_63_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_63_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_63_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_76_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_76_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_76_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_88_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_88_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_88_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_101_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_101_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_101_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_113_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_113_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_113_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_126_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_126_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_126_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_361_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_361_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_361_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_138_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_138_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_151_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_151_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_151_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_163_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_163_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_163_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_176_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_176_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_176_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_188_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_188_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_188_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_201_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_201_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_201_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_261_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_261_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_261_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_274_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_274_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_274_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_286_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_286_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_286_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_299_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_299_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_299_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_311_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_311_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_311_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_324_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_324_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_324_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_336_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_336_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_336_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_349_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_349_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_349_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_374_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_374_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_374_Update/cr
      -- 
    rr_133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_0); -- 
    cr_152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_38_inst_req_1); -- 
    cr_180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_51_inst_req_1); -- 
    cr_208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_63_inst_req_1); -- 
    cr_236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_76_inst_req_1); -- 
    cr_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_88_inst_req_1); -- 
    cr_292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_101_inst_req_1); -- 
    cr_320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_113_inst_req_1); -- 
    cr_348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_126_inst_req_1); -- 
    cr_768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_361_inst_req_1); -- 
    cr_376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_138_inst_req_1); -- 
    cr_404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_151_inst_req_1); -- 
    cr_432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_163_inst_req_1); -- 
    cr_460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_176_inst_req_1); -- 
    cr_488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_188_inst_req_1); -- 
    cr_516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_201_inst_req_1); -- 
    cr_544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_261_inst_req_1); -- 
    cr_572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_274_inst_req_1); -- 
    cr_600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_286_inst_req_1); -- 
    cr_628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_299_inst_req_1); -- 
    cr_656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_311_inst_req_1); -- 
    cr_684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_324_inst_req_1); -- 
    cr_712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_336_inst_req_1); -- 
    cr_740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_349_inst_req_1); -- 
    cr_796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(0), ack => type_cast_374_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_34_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_34_update_start_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_34_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_34_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_34_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_34_Update/cr
      -- 
    ra_134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_0, ack => convTranspose_CP_39_elements(1)); -- 
    cr_138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(1), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_47_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_47_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_47_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_34_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_34_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_34_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_38_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_38_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_38_Sample/rr
      -- 
    ca_139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_1, ack => convTranspose_CP_39_elements(2)); -- 
    rr_147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => type_cast_38_inst_req_0); -- 
    rr_161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(2), ack => RPIPE_ConvTranspose_input_pipe_47_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_38_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_38_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_38_Sample/ra
      -- 
    ra_148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_0, ack => convTranspose_CP_39_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	97 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_38_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_38_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_38_Update/ca
      -- 
    ca_153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_1, ack => convTranspose_CP_39_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_47_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_47_update_start_
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_47_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_47_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_47_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_47_Update/cr
      -- 
    ra_162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_47_inst_ack_0, ack => convTranspose_CP_39_elements(5)); -- 
    cr_166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(5), ack => RPIPE_ConvTranspose_input_pipe_47_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_47_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_47_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_47_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_51_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_51_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_51_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_59_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_59_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_59_Sample/rr
      -- 
    ca_167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_47_inst_ack_1, ack => convTranspose_CP_39_elements(6)); -- 
    rr_175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => type_cast_51_inst_req_0); -- 
    rr_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(6), ack => RPIPE_ConvTranspose_input_pipe_59_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_51_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_51_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_51_Sample/ra
      -- 
    ra_176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_51_inst_ack_0, ack => convTranspose_CP_39_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	97 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_51_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_51_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_51_Update/ca
      -- 
    ca_181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_51_inst_ack_1, ack => convTranspose_CP_39_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_59_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_59_update_start_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_59_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_59_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_59_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_59_Update/cr
      -- 
    ra_190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_59_inst_ack_0, ack => convTranspose_CP_39_elements(9)); -- 
    cr_194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(9), ack => RPIPE_ConvTranspose_input_pipe_59_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_59_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_59_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_59_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_63_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_63_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_63_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_72_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_72_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_72_Sample/rr
      -- 
    ca_195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_59_inst_ack_1, ack => convTranspose_CP_39_elements(10)); -- 
    rr_203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => type_cast_63_inst_req_0); -- 
    rr_217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(10), ack => RPIPE_ConvTranspose_input_pipe_72_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_63_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_63_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_63_Sample/ra
      -- 
    ra_204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_0, ack => convTranspose_CP_39_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	97 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_63_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_63_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_63_Update/ca
      -- 
    ca_209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_1, ack => convTranspose_CP_39_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_72_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_72_update_start_
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_72_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_72_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_72_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_72_Update/cr
      -- 
    ra_218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_72_inst_ack_0, ack => convTranspose_CP_39_elements(13)); -- 
    cr_222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(13), ack => RPIPE_ConvTranspose_input_pipe_72_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_72_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_72_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_72_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_76_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_76_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_76_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_84_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_84_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_84_Sample/rr
      -- 
    ca_223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_72_inst_ack_1, ack => convTranspose_CP_39_elements(14)); -- 
    rr_245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => RPIPE_ConvTranspose_input_pipe_84_inst_req_0); -- 
    rr_231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(14), ack => type_cast_76_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_76_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_76_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_76_Sample/ra
      -- 
    ra_232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_0, ack => convTranspose_CP_39_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	97 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_76_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_76_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_76_Update/ca
      -- 
    ca_237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_1, ack => convTranspose_CP_39_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_84_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_84_update_start_
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_84_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_84_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_84_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_84_Update/cr
      -- 
    ra_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_84_inst_ack_0, ack => convTranspose_CP_39_elements(17)); -- 
    cr_250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(17), ack => RPIPE_ConvTranspose_input_pipe_84_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_84_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_84_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_84_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_88_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_88_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_88_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_97_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_97_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_97_Sample/rr
      -- 
    ca_251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_84_inst_ack_1, ack => convTranspose_CP_39_elements(18)); -- 
    rr_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => type_cast_88_inst_req_0); -- 
    rr_273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(18), ack => RPIPE_ConvTranspose_input_pipe_97_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_88_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_88_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_88_Sample/ra
      -- 
    ra_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_88_inst_ack_0, ack => convTranspose_CP_39_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	97 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_88_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_88_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_88_Update/ca
      -- 
    ca_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_88_inst_ack_1, ack => convTranspose_CP_39_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_97_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_97_update_start_
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_97_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_97_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_97_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_97_Update/cr
      -- 
    ra_274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_97_inst_ack_0, ack => convTranspose_CP_39_elements(21)); -- 
    cr_278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(21), ack => RPIPE_ConvTranspose_input_pipe_97_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_97_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_97_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_97_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_101_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_101_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_101_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_109_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_109_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_109_Sample/rr
      -- 
    ca_279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_97_inst_ack_1, ack => convTranspose_CP_39_elements(22)); -- 
    rr_301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => RPIPE_ConvTranspose_input_pipe_109_inst_req_0); -- 
    rr_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(22), ack => type_cast_101_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_101_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_101_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_101_Sample/ra
      -- 
    ra_288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_101_inst_ack_0, ack => convTranspose_CP_39_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	97 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_101_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_101_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_101_Update/ca
      -- 
    ca_293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_101_inst_ack_1, ack => convTranspose_CP_39_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_109_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_109_update_start_
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_109_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_109_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_109_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_109_Update/cr
      -- 
    ra_302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_109_inst_ack_0, ack => convTranspose_CP_39_elements(25)); -- 
    cr_306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(25), ack => RPIPE_ConvTranspose_input_pipe_109_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_109_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_109_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_109_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_113_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_113_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_113_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_122_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_122_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_122_Sample/rr
      -- 
    ca_307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_109_inst_ack_1, ack => convTranspose_CP_39_elements(26)); -- 
    rr_315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => type_cast_113_inst_req_0); -- 
    rr_329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(26), ack => RPIPE_ConvTranspose_input_pipe_122_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_113_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_113_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_113_Sample/ra
      -- 
    ra_316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_113_inst_ack_0, ack => convTranspose_CP_39_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	97 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_113_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_113_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_113_Update/ca
      -- 
    ca_321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_113_inst_ack_1, ack => convTranspose_CP_39_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_122_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_122_update_start_
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_122_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_122_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_122_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_122_Update/cr
      -- 
    ra_330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_122_inst_ack_0, ack => convTranspose_CP_39_elements(29)); -- 
    cr_334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(29), ack => RPIPE_ConvTranspose_input_pipe_122_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	33 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_134_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_122_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_122_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_122_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_126_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_126_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_126_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_134_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_134_Sample/$entry
      -- 
    ca_335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_122_inst_ack_1, ack => convTranspose_CP_39_elements(30)); -- 
    rr_343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => type_cast_126_inst_req_0); -- 
    rr_357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(30), ack => RPIPE_ConvTranspose_input_pipe_134_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_126_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_126_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_126_Sample/ra
      -- 
    ra_344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_0, ack => convTranspose_CP_39_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	97 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_126_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_126_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_126_Update/ca
      -- 
    ca_349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_126_inst_ack_1, ack => convTranspose_CP_39_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_134_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_134_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_134_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_134_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_134_update_start_
      -- CP-element group 33: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_134_Sample/$exit
      -- 
    ra_358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_134_inst_ack_0, ack => convTranspose_CP_39_elements(33)); -- 
    cr_362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(33), ack => RPIPE_ConvTranspose_input_pipe_134_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_134_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_134_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_138_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_134_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_138_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_138_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_147_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_147_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_147_Sample/rr
      -- 
    ca_363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_134_inst_ack_1, ack => convTranspose_CP_39_elements(34)); -- 
    rr_371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => type_cast_138_inst_req_0); -- 
    rr_385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(34), ack => RPIPE_ConvTranspose_input_pipe_147_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_138_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_138_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_138_Sample/ra
      -- 
    ra_372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_138_inst_ack_0, ack => convTranspose_CP_39_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	97 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_138_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_138_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_138_Update/ca
      -- 
    ca_377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_138_inst_ack_1, ack => convTranspose_CP_39_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_147_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_147_update_start_
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_147_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_147_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_147_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_147_Update/cr
      -- 
    ra_386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_147_inst_ack_0, ack => convTranspose_CP_39_elements(37)); -- 
    cr_390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(37), ack => RPIPE_ConvTranspose_input_pipe_147_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_147_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_147_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_147_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_151_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_151_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_151_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_159_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_159_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_159_Sample/rr
      -- 
    ca_391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_147_inst_ack_1, ack => convTranspose_CP_39_elements(38)); -- 
    rr_399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => type_cast_151_inst_req_0); -- 
    rr_413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(38), ack => RPIPE_ConvTranspose_input_pipe_159_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_151_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_151_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_151_Sample/ra
      -- 
    ra_400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_151_inst_ack_0, ack => convTranspose_CP_39_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	97 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_151_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_151_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_151_Update/ca
      -- 
    ca_405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_151_inst_ack_1, ack => convTranspose_CP_39_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_159_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_159_update_start_
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_159_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_159_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_159_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_159_Update/cr
      -- 
    ra_414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_159_inst_ack_0, ack => convTranspose_CP_39_elements(41)); -- 
    cr_418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(41), ack => RPIPE_ConvTranspose_input_pipe_159_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_159_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_159_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_159_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_163_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_163_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_163_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_172_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_172_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_172_Sample/rr
      -- 
    ca_419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_159_inst_ack_1, ack => convTranspose_CP_39_elements(42)); -- 
    rr_427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => type_cast_163_inst_req_0); -- 
    rr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(42), ack => RPIPE_ConvTranspose_input_pipe_172_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_163_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_163_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_163_Sample/ra
      -- 
    ra_428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_163_inst_ack_0, ack => convTranspose_CP_39_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	97 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_163_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_163_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_163_Update/ca
      -- 
    ca_433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_163_inst_ack_1, ack => convTranspose_CP_39_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_172_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_172_update_start_
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_172_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_172_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_172_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_172_Update/cr
      -- 
    ra_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_172_inst_ack_0, ack => convTranspose_CP_39_elements(45)); -- 
    cr_446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(45), ack => RPIPE_ConvTranspose_input_pipe_172_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_172_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_172_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_172_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_176_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_176_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_176_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_184_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_184_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_184_Sample/rr
      -- 
    ca_447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_172_inst_ack_1, ack => convTranspose_CP_39_elements(46)); -- 
    rr_455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => type_cast_176_inst_req_0); -- 
    rr_469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(46), ack => RPIPE_ConvTranspose_input_pipe_184_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_176_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_176_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_176_Sample/ra
      -- 
    ra_456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_176_inst_ack_0, ack => convTranspose_CP_39_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	97 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_176_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_176_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_176_Update/ca
      -- 
    ca_461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_176_inst_ack_1, ack => convTranspose_CP_39_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_184_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_184_update_start_
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_184_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_184_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_184_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_184_Update/cr
      -- 
    ra_470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_184_inst_ack_0, ack => convTranspose_CP_39_elements(49)); -- 
    cr_474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(49), ack => RPIPE_ConvTranspose_input_pipe_184_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_184_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_184_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_184_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_188_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_188_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_188_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_197_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_197_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_197_Sample/rr
      -- 
    ca_475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_184_inst_ack_1, ack => convTranspose_CP_39_elements(50)); -- 
    rr_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => type_cast_188_inst_req_0); -- 
    rr_497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(50), ack => RPIPE_ConvTranspose_input_pipe_197_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_188_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_188_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_188_Sample/ra
      -- 
    ra_484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_188_inst_ack_0, ack => convTranspose_CP_39_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	97 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_188_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_188_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_188_Update/ca
      -- 
    ca_489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_188_inst_ack_1, ack => convTranspose_CP_39_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_197_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_197_update_start_
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_197_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_197_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_197_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_197_Update/cr
      -- 
    ra_498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_197_inst_ack_0, ack => convTranspose_CP_39_elements(53)); -- 
    cr_502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(53), ack => RPIPE_ConvTranspose_input_pipe_197_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	57 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_197_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_197_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_197_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_201_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_201_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_201_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_257_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_257_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_257_Sample/rr
      -- 
    ca_503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_197_inst_ack_1, ack => convTranspose_CP_39_elements(54)); -- 
    rr_511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => type_cast_201_inst_req_0); -- 
    rr_525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(54), ack => RPIPE_ConvTranspose_input_pipe_257_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_201_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_201_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_201_Sample/ra
      -- 
    ra_512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_201_inst_ack_0, ack => convTranspose_CP_39_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	97 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_201_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_201_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_201_Update/ca
      -- 
    ca_517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_201_inst_ack_1, ack => convTranspose_CP_39_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_257_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_257_update_start_
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_257_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_257_Sample/ra
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_257_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_257_Update/cr
      -- 
    ra_526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_257_inst_ack_0, ack => convTranspose_CP_39_elements(57)); -- 
    cr_530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(57), ack => RPIPE_ConvTranspose_input_pipe_257_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	61 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_257_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_257_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_257_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_261_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_261_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_261_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_270_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_270_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_270_Sample/rr
      -- 
    ca_531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_257_inst_ack_1, ack => convTranspose_CP_39_elements(58)); -- 
    rr_539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(58), ack => type_cast_261_inst_req_0); -- 
    rr_553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(58), ack => RPIPE_ConvTranspose_input_pipe_270_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_261_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_261_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_261_Sample/ra
      -- 
    ra_540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_261_inst_ack_0, ack => convTranspose_CP_39_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	97 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_261_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_261_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_261_Update/ca
      -- 
    ca_545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_261_inst_ack_1, ack => convTranspose_CP_39_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	58 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_270_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_270_update_start_
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_270_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_270_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_270_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_270_Update/cr
      -- 
    ra_554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_270_inst_ack_0, ack => convTranspose_CP_39_elements(61)); -- 
    cr_558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(61), ack => RPIPE_ConvTranspose_input_pipe_270_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	65 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (9) 
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_270_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_270_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_270_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_274_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_274_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_274_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_282_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_282_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_282_Sample/rr
      -- 
    ca_559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_270_inst_ack_1, ack => convTranspose_CP_39_elements(62)); -- 
    rr_581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(62), ack => RPIPE_ConvTranspose_input_pipe_282_inst_req_0); -- 
    rr_567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(62), ack => type_cast_274_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_274_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_274_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_274_Sample/ra
      -- 
    ra_568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_274_inst_ack_0, ack => convTranspose_CP_39_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	0 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	97 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_274_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_274_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_274_Update/ca
      -- 
    ca_573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_274_inst_ack_1, ack => convTranspose_CP_39_elements(64)); -- 
    -- CP-element group 65:  transition  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	62 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (6) 
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_282_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_282_update_start_
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_282_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_282_Sample/ra
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_282_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_282_Update/cr
      -- 
    ra_582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_282_inst_ack_0, ack => convTranspose_CP_39_elements(65)); -- 
    cr_586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(65), ack => RPIPE_ConvTranspose_input_pipe_282_inst_req_1); -- 
    -- CP-element group 66:  fork  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: 	69 
    -- CP-element group 66:  members (9) 
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_282_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_282_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_282_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_286_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_286_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_286_Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_295_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_295_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_295_Sample/rr
      -- 
    ca_587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_282_inst_ack_1, ack => convTranspose_CP_39_elements(66)); -- 
    rr_595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(66), ack => type_cast_286_inst_req_0); -- 
    rr_609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(66), ack => RPIPE_ConvTranspose_input_pipe_295_inst_req_0); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_286_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_286_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_286_Sample/ra
      -- 
    ra_596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_286_inst_ack_0, ack => convTranspose_CP_39_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	97 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_286_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_286_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_286_Update/ca
      -- 
    ca_601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_286_inst_ack_1, ack => convTranspose_CP_39_elements(68)); -- 
    -- CP-element group 69:  transition  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	66 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (6) 
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_295_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_295_update_start_
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_295_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_295_Sample/ra
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_295_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_295_Update/cr
      -- 
    ra_610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_295_inst_ack_0, ack => convTranspose_CP_39_elements(69)); -- 
    cr_614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(69), ack => RPIPE_ConvTranspose_input_pipe_295_inst_req_1); -- 
    -- CP-element group 70:  fork  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	73 
    -- CP-element group 70:  members (9) 
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_295_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_295_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_295_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_299_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_299_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_299_Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_307_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_307_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_307_Sample/rr
      -- 
    ca_615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_295_inst_ack_1, ack => convTranspose_CP_39_elements(70)); -- 
    rr_623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(70), ack => type_cast_299_inst_req_0); -- 
    rr_637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(70), ack => RPIPE_ConvTranspose_input_pipe_307_inst_req_0); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_299_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_299_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_299_Sample/ra
      -- 
    ra_624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_299_inst_ack_0, ack => convTranspose_CP_39_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	0 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	97 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_299_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_299_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_299_Update/ca
      -- 
    ca_629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_299_inst_ack_1, ack => convTranspose_CP_39_elements(72)); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	70 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_307_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_307_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_307_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_307_Sample/ra
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_307_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_307_Update/cr
      -- 
    ra_638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_307_inst_ack_0, ack => convTranspose_CP_39_elements(73)); -- 
    cr_642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(73), ack => RPIPE_ConvTranspose_input_pipe_307_inst_req_1); -- 
    -- CP-element group 74:  fork  transition  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	77 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (9) 
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_307_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_307_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_307_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_311_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_311_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_311_Sample/rr
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_320_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_320_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_320_Sample/rr
      -- 
    ca_643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_307_inst_ack_1, ack => convTranspose_CP_39_elements(74)); -- 
    rr_651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(74), ack => type_cast_311_inst_req_0); -- 
    rr_665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(74), ack => RPIPE_ConvTranspose_input_pipe_320_inst_req_0); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_311_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_311_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_311_Sample/ra
      -- 
    ra_652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_311_inst_ack_0, ack => convTranspose_CP_39_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	0 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	97 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_311_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_311_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_311_Update/ca
      -- 
    ca_657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_311_inst_ack_1, ack => convTranspose_CP_39_elements(76)); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	74 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_320_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_320_update_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_320_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_320_Sample/ra
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_320_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_320_Update/cr
      -- 
    ra_666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_320_inst_ack_0, ack => convTranspose_CP_39_elements(77)); -- 
    cr_670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(77), ack => RPIPE_ConvTranspose_input_pipe_320_inst_req_1); -- 
    -- CP-element group 78:  fork  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	81 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (9) 
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_320_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_320_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_320_Update/ca
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_324_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_324_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_324_Sample/rr
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_332_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_332_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_332_Sample/rr
      -- 
    ca_671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_320_inst_ack_1, ack => convTranspose_CP_39_elements(78)); -- 
    rr_679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(78), ack => type_cast_324_inst_req_0); -- 
    rr_693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(78), ack => RPIPE_ConvTranspose_input_pipe_332_inst_req_0); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_324_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_324_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_324_Sample/ra
      -- 
    ra_680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_324_inst_ack_0, ack => convTranspose_CP_39_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	0 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	97 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_324_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_324_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_324_Update/ca
      -- 
    ca_685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_324_inst_ack_1, ack => convTranspose_CP_39_elements(80)); -- 
    -- CP-element group 81:  transition  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	78 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (6) 
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_332_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_332_update_start_
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_332_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_332_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_332_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_332_Update/cr
      -- 
    ra_694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_332_inst_ack_0, ack => convTranspose_CP_39_elements(81)); -- 
    cr_698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(81), ack => RPIPE_ConvTranspose_input_pipe_332_inst_req_1); -- 
    -- CP-element group 82:  fork  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82: 	85 
    -- CP-element group 82:  members (9) 
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_332_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_332_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_332_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_336_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_336_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_336_Sample/rr
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_345_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_345_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_345_Sample/rr
      -- 
    ca_699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_332_inst_ack_1, ack => convTranspose_CP_39_elements(82)); -- 
    rr_707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(82), ack => type_cast_336_inst_req_0); -- 
    rr_721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(82), ack => RPIPE_ConvTranspose_input_pipe_345_inst_req_0); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_336_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_336_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_336_Sample/ra
      -- 
    ra_708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_336_inst_ack_0, ack => convTranspose_CP_39_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	0 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	97 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_336_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_336_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_336_Update/ca
      -- 
    ca_713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_336_inst_ack_1, ack => convTranspose_CP_39_elements(84)); -- 
    -- CP-element group 85:  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	82 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_345_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_345_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_345_update_start_
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_345_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_345_Sample/ra
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_345_Update/cr
      -- 
    ra_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_345_inst_ack_0, ack => convTranspose_CP_39_elements(85)); -- 
    cr_726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(85), ack => RPIPE_ConvTranspose_input_pipe_345_inst_req_1); -- 
    -- CP-element group 86:  fork  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86: 	89 
    -- CP-element group 86:  members (9) 
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_345_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_345_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_345_Update/ca
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_349_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_349_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_349_Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_357_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_357_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_357_Sample/rr
      -- 
    ca_727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_345_inst_ack_1, ack => convTranspose_CP_39_elements(86)); -- 
    rr_735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(86), ack => type_cast_349_inst_req_0); -- 
    rr_749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(86), ack => RPIPE_ConvTranspose_input_pipe_357_inst_req_0); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_349_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_349_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_349_Sample/ra
      -- 
    ra_736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_349_inst_ack_0, ack => convTranspose_CP_39_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	0 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	97 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_349_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_349_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_349_Update/ca
      -- 
    ca_741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_349_inst_ack_1, ack => convTranspose_CP_39_elements(88)); -- 
    -- CP-element group 89:  transition  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	86 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89:  members (6) 
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_357_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_357_update_start_
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_357_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_357_Sample/ra
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_357_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_357_Update/cr
      -- 
    ra_750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_357_inst_ack_0, ack => convTranspose_CP_39_elements(89)); -- 
    cr_754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(89), ack => RPIPE_ConvTranspose_input_pipe_357_inst_req_1); -- 
    -- CP-element group 90:  fork  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90: 	93 
    -- CP-element group 90:  members (9) 
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_361_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_361_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_361_Sample/rr
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_370_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_370_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_370_Sample/rr
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_357_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_357_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_357_Update/ca
      -- 
    ca_755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_357_inst_ack_1, ack => convTranspose_CP_39_elements(90)); -- 
    rr_763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(90), ack => type_cast_361_inst_req_0); -- 
    rr_777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(90), ack => RPIPE_ConvTranspose_input_pipe_370_inst_req_0); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_361_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_361_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_361_Sample/ra
      -- 
    ra_764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_361_inst_ack_0, ack => convTranspose_CP_39_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	0 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	97 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_361_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_361_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_361_Update/ca
      -- 
    ca_769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_361_inst_ack_1, ack => convTranspose_CP_39_elements(92)); -- 
    -- CP-element group 93:  transition  input  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	90 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (6) 
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_370_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_370_update_start_
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_370_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_370_Sample/ra
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_370_Update/$entry
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_370_Update/cr
      -- 
    ra_778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_370_inst_ack_0, ack => convTranspose_CP_39_elements(93)); -- 
    cr_782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(93), ack => RPIPE_ConvTranspose_input_pipe_370_inst_req_1); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_370_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_370_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/RPIPE_ConvTranspose_input_pipe_370_Update/ca
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_374_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_374_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_374_Sample/rr
      -- 
    ca_783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_370_inst_ack_1, ack => convTranspose_CP_39_elements(94)); -- 
    rr_791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(94), ack => type_cast_374_inst_req_0); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_374_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_374_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_374_Sample/ra
      -- 
    ra_792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_374_inst_ack_0, ack => convTranspose_CP_39_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	0 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_374_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_374_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/type_cast_374_Update/ca
      -- 
    ca_797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_374_inst_ack_1, ack => convTranspose_CP_39_elements(96)); -- 
    -- CP-element group 97:  branch  join  transition  place  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	24 
    -- CP-element group 97: 	20 
    -- CP-element group 97: 	32 
    -- CP-element group 97: 	28 
    -- CP-element group 97: 	16 
    -- CP-element group 97: 	84 
    -- CP-element group 97: 	88 
    -- CP-element group 97: 	80 
    -- CP-element group 97: 	92 
    -- CP-element group 97: 	96 
    -- CP-element group 97: 	68 
    -- CP-element group 97: 	72 
    -- CP-element group 97: 	76 
    -- CP-element group 97: 	36 
    -- CP-element group 97: 	40 
    -- CP-element group 97: 	44 
    -- CP-element group 97: 	48 
    -- CP-element group 97: 	52 
    -- CP-element group 97: 	56 
    -- CP-element group 97: 	60 
    -- CP-element group 97: 	64 
    -- CP-element group 97: 	4 
    -- CP-element group 97: 	8 
    -- CP-element group 97: 	12 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (10) 
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387__exit__
      -- CP-element group 97: 	 branch_block_stmt_32/if_stmt_388__entry__
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_387/$exit
      -- CP-element group 97: 	 branch_block_stmt_32/if_stmt_388_dead_link/$entry
      -- CP-element group 97: 	 branch_block_stmt_32/if_stmt_388_eval_test/$entry
      -- CP-element group 97: 	 branch_block_stmt_32/if_stmt_388_eval_test/$exit
      -- CP-element group 97: 	 branch_block_stmt_32/if_stmt_388_eval_test/branch_req
      -- CP-element group 97: 	 branch_block_stmt_32/R_cmp487_389_place
      -- CP-element group 97: 	 branch_block_stmt_32/if_stmt_388_if_link/$entry
      -- CP-element group 97: 	 branch_block_stmt_32/if_stmt_388_else_link/$entry
      -- 
    branch_req_805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(97), ack => if_stmt_388_branch_req_0); -- 
    convTranspose_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 23) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1);
      constant place_markings: IntegerArray(0 to 23)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0);
      constant place_delays: IntegerArray(0 to 23) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 24); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(24) & convTranspose_CP_39_elements(20) & convTranspose_CP_39_elements(32) & convTranspose_CP_39_elements(28) & convTranspose_CP_39_elements(16) & convTranspose_CP_39_elements(84) & convTranspose_CP_39_elements(88) & convTranspose_CP_39_elements(80) & convTranspose_CP_39_elements(92) & convTranspose_CP_39_elements(96) & convTranspose_CP_39_elements(68) & convTranspose_CP_39_elements(72) & convTranspose_CP_39_elements(76) & convTranspose_CP_39_elements(36) & convTranspose_CP_39_elements(40) & convTranspose_CP_39_elements(44) & convTranspose_CP_39_elements(48) & convTranspose_CP_39_elements(52) & convTranspose_CP_39_elements(56) & convTranspose_CP_39_elements(60) & convTranspose_CP_39_elements(64) & convTranspose_CP_39_elements(4) & convTranspose_CP_39_elements(8) & convTranspose_CP_39_elements(12);
      gj_convTranspose_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 24, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	102 
    -- CP-element group 98: 	103 
    -- CP-element group 98:  members (18) 
      -- CP-element group 98: 	 branch_block_stmt_32/merge_stmt_409__exit__
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_415_to_assign_stmt_438__entry__
      -- CP-element group 98: 	 branch_block_stmt_32/merge_stmt_409_PhiReqMerge
      -- CP-element group 98: 	 branch_block_stmt_32/if_stmt_388_if_link/$exit
      -- CP-element group 98: 	 branch_block_stmt_32/if_stmt_388_if_link/if_choice_transition
      -- CP-element group 98: 	 branch_block_stmt_32/entry_bbx_xnph489
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_415_to_assign_stmt_438/$entry
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_415_to_assign_stmt_438/type_cast_424_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_415_to_assign_stmt_438/type_cast_424_update_start_
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_415_to_assign_stmt_438/type_cast_424_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_415_to_assign_stmt_438/type_cast_424_Sample/rr
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_415_to_assign_stmt_438/type_cast_424_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_415_to_assign_stmt_438/type_cast_424_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_32/merge_stmt_409_PhiAck/dummy
      -- CP-element group 98: 	 branch_block_stmt_32/merge_stmt_409_PhiAck/$exit
      -- CP-element group 98: 	 branch_block_stmt_32/merge_stmt_409_PhiAck/$entry
      -- CP-element group 98: 	 branch_block_stmt_32/entry_bbx_xnph489_PhiReq/$exit
      -- CP-element group 98: 	 branch_block_stmt_32/entry_bbx_xnph489_PhiReq/$entry
      -- 
    if_choice_transition_810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_388_branch_ack_1, ack => convTranspose_CP_39_elements(98)); -- 
    rr_849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(98), ack => type_cast_424_inst_req_0); -- 
    cr_854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(98), ack => type_cast_424_inst_req_1); -- 
    -- CP-element group 99:  transition  place  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	378 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_32/if_stmt_388_else_link/$exit
      -- CP-element group 99: 	 branch_block_stmt_32/if_stmt_388_else_link/else_choice_transition
      -- CP-element group 99: 	 branch_block_stmt_32/entry_forx_xcond190x_xpreheader
      -- CP-element group 99: 	 branch_block_stmt_32/entry_forx_xcond190x_xpreheader_PhiReq/$exit
      -- CP-element group 99: 	 branch_block_stmt_32/entry_forx_xcond190x_xpreheader_PhiReq/$entry
      -- 
    else_choice_transition_814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_388_branch_ack_0, ack => convTranspose_CP_39_elements(99)); -- 
    -- CP-element group 100:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	378 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	146 
    -- CP-element group 100: 	147 
    -- CP-element group 100:  members (18) 
      -- CP-element group 100: 	 branch_block_stmt_32/merge_stmt_610__exit__
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_616_to_assign_stmt_645__entry__
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_616_to_assign_stmt_645/type_cast_631_update_start_
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_616_to_assign_stmt_645/type_cast_631_Update/cr
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_616_to_assign_stmt_645/type_cast_631_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_616_to_assign_stmt_645/type_cast_631_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_616_to_assign_stmt_645/type_cast_631_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_616_to_assign_stmt_645/type_cast_631_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_616_to_assign_stmt_645/$entry
      -- CP-element group 100: 	 branch_block_stmt_32/if_stmt_403_if_link/$exit
      -- CP-element group 100: 	 branch_block_stmt_32/if_stmt_403_if_link/if_choice_transition
      -- CP-element group 100: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_bbx_xnph485
      -- CP-element group 100: 	 branch_block_stmt_32/merge_stmt_610_PhiReqMerge
      -- CP-element group 100: 	 branch_block_stmt_32/merge_stmt_610_PhiAck/dummy
      -- CP-element group 100: 	 branch_block_stmt_32/merge_stmt_610_PhiAck/$exit
      -- CP-element group 100: 	 branch_block_stmt_32/merge_stmt_610_PhiAck/$entry
      -- CP-element group 100: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_bbx_xnph485_PhiReq/$exit
      -- CP-element group 100: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_bbx_xnph485_PhiReq/$entry
      -- 
    if_choice_transition_832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_403_branch_ack_1, ack => convTranspose_CP_39_elements(100)); -- 
    cr_1213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(100), ack => type_cast_631_inst_req_1); -- 
    rr_1208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(100), ack => type_cast_631_inst_req_0); -- 
    -- CP-element group 101:  transition  place  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	378 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	391 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$entry
      -- CP-element group 101: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_forx_xend250_PhiReq/$exit
      -- CP-element group 101: 	 branch_block_stmt_32/if_stmt_403_else_link/$exit
      -- CP-element group 101: 	 branch_block_stmt_32/if_stmt_403_else_link/else_choice_transition
      -- CP-element group 101: 	 branch_block_stmt_32/forx_xcond190x_xpreheader_forx_xend250
      -- 
    else_choice_transition_836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_403_branch_ack_0, ack => convTranspose_CP_39_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	98 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_415_to_assign_stmt_438/type_cast_424_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_415_to_assign_stmt_438/type_cast_424_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_415_to_assign_stmt_438/type_cast_424_Sample/ra
      -- 
    ra_850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_424_inst_ack_0, ack => convTranspose_CP_39_elements(102)); -- 
    -- CP-element group 103:  transition  place  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	98 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	379 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_415_to_assign_stmt_438__exit__
      -- CP-element group 103: 	 branch_block_stmt_32/bbx_xnph489_forx_xbody
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_415_to_assign_stmt_438/$exit
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_415_to_assign_stmt_438/type_cast_424_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_415_to_assign_stmt_438/type_cast_424_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_415_to_assign_stmt_438/type_cast_424_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_32/bbx_xnph489_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/$entry
      -- CP-element group 103: 	 branch_block_stmt_32/bbx_xnph489_forx_xbody_PhiReq/phi_stmt_441/$entry
      -- CP-element group 103: 	 branch_block_stmt_32/bbx_xnph489_forx_xbody_PhiReq/$entry
      -- 
    ca_855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_424_inst_ack_1, ack => convTranspose_CP_39_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	384 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	143 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_final_index_sum_regn_sample_complete
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_final_index_sum_regn_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_final_index_sum_regn_Sample/ack
      -- 
    ack_884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_453_index_offset_ack_0, ack => convTranspose_CP_39_elements(104)); -- 
    -- CP-element group 105:  transition  input  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	384 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (11) 
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/addr_of_454_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_root_address_calculated
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_offset_calculated
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_final_index_sum_regn_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_final_index_sum_regn_Update/ack
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_base_plus_offset/$entry
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_base_plus_offset/$exit
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_base_plus_offset/sum_rename_req
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_base_plus_offset/sum_rename_ack
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/addr_of_454_request/$entry
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/addr_of_454_request/req
      -- 
    ack_889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_453_index_offset_ack_1, ack => convTranspose_CP_39_elements(105)); -- 
    req_898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(105), ack => addr_of_454_final_reg_req_0); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/addr_of_454_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/addr_of_454_request/$exit
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/addr_of_454_request/ack
      -- 
    ack_899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_454_final_reg_ack_0, ack => convTranspose_CP_39_elements(106)); -- 
    -- CP-element group 107:  fork  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	384 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	140 
    -- CP-element group 107:  members (19) 
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_base_address_resized
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_root_address_calculated
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_word_addrgen/root_register_ack
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_word_addrgen/root_register_req
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_word_addrgen/$exit
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_word_addrgen/$entry
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_base_plus_offset/sum_rename_ack
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_base_plus_offset/sum_rename_req
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_base_plus_offset/$exit
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_base_plus_offset/$entry
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_base_addr_resize/base_resize_ack
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_base_addr_resize/base_resize_req
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_base_addr_resize/$exit
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_base_addr_resize/$entry
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_word_address_calculated
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_base_address_calculated
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/addr_of_454_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/addr_of_454_complete/$exit
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/addr_of_454_complete/ack
      -- 
    ack_904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_454_final_reg_ack_1, ack => convTranspose_CP_39_elements(107)); -- 
    -- CP-element group 108:  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	384 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (6) 
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_457_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_457_update_start_
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_457_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_457_Sample/ra
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_457_Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_457_Update/cr
      -- 
    ra_913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_457_inst_ack_0, ack => convTranspose_CP_39_elements(108)); -- 
    cr_917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(108), ack => RPIPE_ConvTranspose_input_pipe_457_inst_req_1); -- 
    -- CP-element group 109:  fork  transition  input  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109: 	112 
    -- CP-element group 109:  members (9) 
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_457_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_457_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_457_Update/ca
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_461_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_461_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_461_Sample/rr
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_470_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_470_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_470_Sample/rr
      -- 
    ca_918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_457_inst_ack_1, ack => convTranspose_CP_39_elements(109)); -- 
    rr_926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(109), ack => type_cast_461_inst_req_0); -- 
    rr_940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(109), ack => RPIPE_ConvTranspose_input_pipe_470_inst_req_0); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_461_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_461_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_461_Sample/ra
      -- 
    ra_927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_461_inst_ack_0, ack => convTranspose_CP_39_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	384 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	140 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_461_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_461_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_461_Update/ca
      -- 
    ca_932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_461_inst_ack_1, ack => convTranspose_CP_39_elements(111)); -- 
    -- CP-element group 112:  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	109 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (6) 
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_470_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_470_update_start_
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_470_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_470_Sample/ra
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_470_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_470_Update/cr
      -- 
    ra_941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_470_inst_ack_0, ack => convTranspose_CP_39_elements(112)); -- 
    cr_945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(112), ack => RPIPE_ConvTranspose_input_pipe_470_inst_req_1); -- 
    -- CP-element group 113:  fork  transition  input  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	116 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (9) 
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_488_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_488_Sample/rr
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_488_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_470_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_470_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_470_Update/ca
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_474_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_474_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_474_Sample/rr
      -- 
    ca_946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_470_inst_ack_1, ack => convTranspose_CP_39_elements(113)); -- 
    rr_968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(113), ack => RPIPE_ConvTranspose_input_pipe_488_inst_req_0); -- 
    rr_954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(113), ack => type_cast_474_inst_req_0); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_474_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_474_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_474_Sample/ra
      -- 
    ra_955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_474_inst_ack_0, ack => convTranspose_CP_39_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	384 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	140 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_474_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_474_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_474_update_completed_
      -- 
    ca_960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_474_inst_ack_1, ack => convTranspose_CP_39_elements(115)); -- 
    -- CP-element group 116:  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	113 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (6) 
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_488_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_488_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_488_Sample/ra
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_488_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_488_update_start_
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_488_sample_completed_
      -- 
    ra_969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_488_inst_ack_0, ack => convTranspose_CP_39_elements(116)); -- 
    cr_973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(116), ack => RPIPE_ConvTranspose_input_pipe_488_inst_req_1); -- 
    -- CP-element group 117:  fork  transition  input  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117: 	120 
    -- CP-element group 117:  members (9) 
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_492_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_488_Update/ca
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_488_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_488_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_506_Sample/rr
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_506_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_506_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_492_Sample/rr
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_492_Sample/$entry
      -- 
    ca_974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_488_inst_ack_1, ack => convTranspose_CP_39_elements(117)); -- 
    rr_982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(117), ack => type_cast_492_inst_req_0); -- 
    rr_996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(117), ack => RPIPE_ConvTranspose_input_pipe_506_inst_req_0); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_492_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_492_Sample/ra
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_492_Sample/$exit
      -- 
    ra_983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_492_inst_ack_0, ack => convTranspose_CP_39_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	384 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	140 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_492_Update/ca
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_492_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_492_update_completed_
      -- 
    ca_988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_492_inst_ack_1, ack => convTranspose_CP_39_elements(119)); -- 
    -- CP-element group 120:  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	117 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (6) 
      -- CP-element group 120: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_506_Update/cr
      -- CP-element group 120: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_506_Update/$entry
      -- CP-element group 120: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_506_Sample/ra
      -- CP-element group 120: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_506_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_506_update_start_
      -- CP-element group 120: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_506_sample_completed_
      -- 
    ra_997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_506_inst_ack_0, ack => convTranspose_CP_39_elements(120)); -- 
    cr_1001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(120), ack => RPIPE_ConvTranspose_input_pipe_506_inst_req_1); -- 
    -- CP-element group 121:  fork  transition  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: 	124 
    -- CP-element group 121:  members (9) 
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_524_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_524_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_524_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_510_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_510_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_510_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_506_Update/ca
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_506_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_506_update_completed_
      -- 
    ca_1002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_506_inst_ack_1, ack => convTranspose_CP_39_elements(121)); -- 
    rr_1010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => type_cast_510_inst_req_0); -- 
    rr_1024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(121), ack => RPIPE_ConvTranspose_input_pipe_524_inst_req_0); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_510_Sample/ra
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_510_Sample/$exit
      -- CP-element group 122: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_510_sample_completed_
      -- 
    ra_1011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_510_inst_ack_0, ack => convTranspose_CP_39_elements(122)); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	384 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	140 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_510_Update/ca
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_510_Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_510_update_completed_
      -- 
    ca_1016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_510_inst_ack_1, ack => convTranspose_CP_39_elements(123)); -- 
    -- CP-element group 124:  transition  input  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (6) 
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_524_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_524_Sample/ra
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_524_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_524_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_524_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_524_update_start_
      -- 
    ra_1025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_524_inst_ack_0, ack => convTranspose_CP_39_elements(124)); -- 
    cr_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(124), ack => RPIPE_ConvTranspose_input_pipe_524_inst_req_1); -- 
    -- CP-element group 125:  fork  transition  input  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125: 	128 
    -- CP-element group 125:  members (9) 
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_528_Sample/rr
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_542_Sample/rr
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_528_Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_542_Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_542_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_528_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_524_Update/ca
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_524_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_524_update_completed_
      -- 
    ca_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_524_inst_ack_1, ack => convTranspose_CP_39_elements(125)); -- 
    rr_1038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(125), ack => type_cast_528_inst_req_0); -- 
    rr_1052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(125), ack => RPIPE_ConvTranspose_input_pipe_542_inst_req_0); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_528_Sample/ra
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_528_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_528_sample_completed_
      -- 
    ra_1039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_528_inst_ack_0, ack => convTranspose_CP_39_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	384 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	140 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_528_Update/ca
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_528_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_528_update_completed_
      -- 
    ca_1044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_528_inst_ack_1, ack => convTranspose_CP_39_elements(127)); -- 
    -- CP-element group 128:  transition  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	125 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (6) 
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_542_Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_542_Sample/ra
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_542_Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_542_update_start_
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_542_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_542_Update/cr
      -- 
    ra_1053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_542_inst_ack_0, ack => convTranspose_CP_39_elements(128)); -- 
    cr_1057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(128), ack => RPIPE_ConvTranspose_input_pipe_542_inst_req_1); -- 
    -- CP-element group 129:  fork  transition  input  output  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129: 	132 
    -- CP-element group 129:  members (9) 
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_542_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_560_Sample/rr
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_560_Sample/$entry
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_560_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_546_Sample/rr
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_546_Sample/$entry
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_546_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_542_Update/ca
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_542_Update/$exit
      -- 
    ca_1058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_542_inst_ack_1, ack => convTranspose_CP_39_elements(129)); -- 
    rr_1066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(129), ack => type_cast_546_inst_req_0); -- 
    rr_1080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(129), ack => RPIPE_ConvTranspose_input_pipe_560_inst_req_0); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_546_Sample/ra
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_546_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_546_sample_completed_
      -- 
    ra_1067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_546_inst_ack_0, ack => convTranspose_CP_39_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	384 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	140 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_546_Update/ca
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_546_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_546_update_completed_
      -- 
    ca_1072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_546_inst_ack_1, ack => convTranspose_CP_39_elements(131)); -- 
    -- CP-element group 132:  transition  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	129 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (6) 
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_560_Update/cr
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_560_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_560_Sample/ra
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_560_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_560_update_start_
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_560_sample_completed_
      -- 
    ra_1081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_560_inst_ack_0, ack => convTranspose_CP_39_elements(132)); -- 
    cr_1085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(132), ack => RPIPE_ConvTranspose_input_pipe_560_inst_req_1); -- 
    -- CP-element group 133:  fork  transition  input  output  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	134 
    -- CP-element group 133: 	136 
    -- CP-element group 133:  members (9) 
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_560_Update/ca
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_560_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_560_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_578_Sample/rr
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_578_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_578_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_564_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_564_Sample/rr
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_564_Sample/$entry
      -- 
    ca_1086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_560_inst_ack_1, ack => convTranspose_CP_39_elements(133)); -- 
    rr_1094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(133), ack => type_cast_564_inst_req_0); -- 
    rr_1108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(133), ack => RPIPE_ConvTranspose_input_pipe_578_inst_req_0); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	133 
    -- CP-element group 134: successors 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_564_Sample/ra
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_564_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_564_Sample/$exit
      -- 
    ra_1095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_564_inst_ack_0, ack => convTranspose_CP_39_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	384 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	140 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_564_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_564_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_564_Update/ca
      -- 
    ca_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_564_inst_ack_1, ack => convTranspose_CP_39_elements(135)); -- 
    -- CP-element group 136:  transition  input  output  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	133 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (6) 
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_578_Update/cr
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_578_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_578_Sample/ra
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_578_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_578_update_start_
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_578_sample_completed_
      -- 
    ra_1109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_578_inst_ack_0, ack => convTranspose_CP_39_elements(136)); -- 
    cr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(136), ack => RPIPE_ConvTranspose_input_pipe_578_inst_req_1); -- 
    -- CP-element group 137:  transition  input  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_582_Sample/rr
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_582_Sample/$entry
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_582_sample_start_
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_578_Update/ca
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_578_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_578_update_completed_
      -- 
    ca_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_578_inst_ack_1, ack => convTranspose_CP_39_elements(137)); -- 
    rr_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(137), ack => type_cast_582_inst_req_0); -- 
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_582_Sample/ra
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_582_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_582_sample_completed_
      -- 
    ra_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_582_inst_ack_0, ack => convTranspose_CP_39_elements(138)); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	384 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_582_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_582_Update/ca
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_582_Update/$exit
      -- 
    ca_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_582_inst_ack_1, ack => convTranspose_CP_39_elements(139)); -- 
    -- CP-element group 140:  join  transition  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	115 
    -- CP-element group 140: 	119 
    -- CP-element group 140: 	123 
    -- CP-element group 140: 	127 
    -- CP-element group 140: 	131 
    -- CP-element group 140: 	135 
    -- CP-element group 140: 	139 
    -- CP-element group 140: 	107 
    -- CP-element group 140: 	111 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	141 
    -- CP-element group 140:  members (9) 
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Sample/ptr_deref_590_Split/split_req
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Sample/ptr_deref_590_Split/$exit
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Sample/word_access_start/word_0/rr
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Sample/word_access_start/word_0/$entry
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Sample/word_access_start/$entry
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Sample/ptr_deref_590_Split/split_ack
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Sample/ptr_deref_590_Split/$entry
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Sample/$entry
      -- 
    rr_1166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(140), ack => ptr_deref_590_store_0_req_0); -- 
    convTranspose_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(115) & convTranspose_CP_39_elements(119) & convTranspose_CP_39_elements(123) & convTranspose_CP_39_elements(127) & convTranspose_CP_39_elements(131) & convTranspose_CP_39_elements(135) & convTranspose_CP_39_elements(139) & convTranspose_CP_39_elements(107) & convTranspose_CP_39_elements(111);
      gj_convTranspose_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	140 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (5) 
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Sample/word_access_start/word_0/ra
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Sample/word_access_start/word_0/$exit
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Sample/word_access_start/$exit
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Sample/$exit
      -- 
    ra_1167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_590_store_0_ack_0, ack => convTranspose_CP_39_elements(141)); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	384 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142:  members (5) 
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Update/word_access_complete/word_0/$exit
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Update/word_access_complete/$exit
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Update/word_access_complete/word_0/ca
      -- 
    ca_1178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_590_store_0_ack_1, ack => convTranspose_CP_39_elements(142)); -- 
    -- CP-element group 143:  branch  join  transition  place  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: 	104 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (10) 
      -- CP-element group 143: 	 branch_block_stmt_32/if_stmt_604_if_link/$entry
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603__exit__
      -- CP-element group 143: 	 branch_block_stmt_32/if_stmt_604__entry__
      -- CP-element group 143: 	 branch_block_stmt_32/R_exitcond3_605_place
      -- CP-element group 143: 	 branch_block_stmt_32/if_stmt_604_eval_test/branch_req
      -- CP-element group 143: 	 branch_block_stmt_32/if_stmt_604_eval_test/$exit
      -- CP-element group 143: 	 branch_block_stmt_32/if_stmt_604_eval_test/$entry
      -- CP-element group 143: 	 branch_block_stmt_32/if_stmt_604_dead_link/$entry
      -- CP-element group 143: 	 branch_block_stmt_32/if_stmt_604_else_link/$entry
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/$exit
      -- 
    branch_req_1186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(143), ack => if_stmt_604_branch_req_0); -- 
    convTranspose_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(142) & convTranspose_CP_39_elements(104);
      gj_convTranspose_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  merge  transition  place  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	378 
    -- CP-element group 144:  members (13) 
      -- CP-element group 144: 	 branch_block_stmt_32/if_stmt_604_if_link/if_choice_transition
      -- CP-element group 144: 	 branch_block_stmt_32/merge_stmt_394_PhiReqMerge
      -- CP-element group 144: 	 branch_block_stmt_32/merge_stmt_394__exit__
      -- CP-element group 144: 	 branch_block_stmt_32/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader
      -- CP-element group 144: 	 branch_block_stmt_32/if_stmt_604_if_link/$exit
      -- CP-element group 144: 	 branch_block_stmt_32/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit
      -- CP-element group 144: 	 branch_block_stmt_32/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$exit
      -- CP-element group 144: 	 branch_block_stmt_32/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 144: 	 branch_block_stmt_32/forx_xcond190x_xpreheaderx_xloopexit_forx_xcond190x_xpreheader_PhiReq/$entry
      -- CP-element group 144: 	 branch_block_stmt_32/merge_stmt_394_PhiAck/dummy
      -- CP-element group 144: 	 branch_block_stmt_32/merge_stmt_394_PhiAck/$exit
      -- CP-element group 144: 	 branch_block_stmt_32/merge_stmt_394_PhiAck/$entry
      -- CP-element group 144: 	 branch_block_stmt_32/forx_xbody_forx_xcond190x_xpreheaderx_xloopexit_PhiReq/$exit
      -- 
    if_choice_transition_1191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_604_branch_ack_1, ack => convTranspose_CP_39_elements(144)); -- 
    -- CP-element group 145:  fork  transition  place  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	380 
    -- CP-element group 145: 	381 
    -- CP-element group 145:  members (12) 
      -- CP-element group 145: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/$entry
      -- CP-element group 145: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/$entry
      -- CP-element group 145: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_32/if_stmt_604_else_link/$exit
      -- CP-element group 145: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/$entry
      -- CP-element group 145: 	 branch_block_stmt_32/if_stmt_604_else_link/else_choice_transition
      -- CP-element group 145: 	 branch_block_stmt_32/forx_xbody_forx_xbody
      -- CP-element group 145: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/$entry
      -- CP-element group 145: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/Sample/rr
      -- CP-element group 145: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 145: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_604_branch_ack_0, ack => convTranspose_CP_39_elements(145)); -- 
    rr_3016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(145), ack => type_cast_447_inst_req_0); -- 
    cr_3021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(145), ack => type_cast_447_inst_req_1); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	100 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_616_to_assign_stmt_645/type_cast_631_Sample/ra
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_616_to_assign_stmt_645/type_cast_631_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_616_to_assign_stmt_645/type_cast_631_sample_completed_
      -- 
    ra_1209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_631_inst_ack_0, ack => convTranspose_CP_39_elements(146)); -- 
    -- CP-element group 147:  transition  place  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	100 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	385 
    -- CP-element group 147:  members (9) 
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_616_to_assign_stmt_645__exit__
      -- CP-element group 147: 	 branch_block_stmt_32/bbx_xnph485_forx_xbody196
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_616_to_assign_stmt_645/type_cast_631_Update/ca
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_616_to_assign_stmt_645/type_cast_631_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_616_to_assign_stmt_645/type_cast_631_update_completed_
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_616_to_assign_stmt_645/$exit
      -- CP-element group 147: 	 branch_block_stmt_32/bbx_xnph485_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_sources/$entry
      -- CP-element group 147: 	 branch_block_stmt_32/bbx_xnph485_forx_xbody196_PhiReq/phi_stmt_648/$entry
      -- CP-element group 147: 	 branch_block_stmt_32/bbx_xnph485_forx_xbody196_PhiReq/$entry
      -- 
    ca_1214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_631_inst_ack_1, ack => convTranspose_CP_39_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	390 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	187 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_final_index_sum_regn_Sample/ack
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_final_index_sum_regn_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_final_index_sum_regn_sample_complete
      -- 
    ack_1243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_660_index_offset_ack_0, ack => convTranspose_CP_39_elements(148)); -- 
    -- CP-element group 149:  transition  input  output  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	390 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (11) 
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_base_plus_offset/sum_rename_ack
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_base_plus_offset/sum_rename_req
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_base_plus_offset/$exit
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_base_plus_offset/$entry
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_offset_calculated
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_root_address_calculated
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_final_index_sum_regn_Update/ack
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_final_index_sum_regn_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/addr_of_661_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/addr_of_661_request/req
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/addr_of_661_request/$entry
      -- 
    ack_1248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_660_index_offset_ack_1, ack => convTranspose_CP_39_elements(149)); -- 
    req_1257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(149), ack => addr_of_661_final_reg_req_0); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/addr_of_661_sample_completed_
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/addr_of_661_request/ack
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/addr_of_661_request/$exit
      -- 
    ack_1258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_661_final_reg_ack_0, ack => convTranspose_CP_39_elements(150)); -- 
    -- CP-element group 151:  fork  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	390 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	184 
    -- CP-element group 151:  members (19) 
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/addr_of_661_update_completed_
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/addr_of_661_complete/ack
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/addr_of_661_complete/$exit
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_base_address_calculated
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_word_address_calculated
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_root_address_calculated
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_base_address_resized
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_base_addr_resize/$entry
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_base_addr_resize/$exit
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_base_addr_resize/base_resize_req
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_base_addr_resize/base_resize_ack
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_base_plus_offset/$entry
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_base_plus_offset/$exit
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_base_plus_offset/sum_rename_req
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_base_plus_offset/sum_rename_ack
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_word_addrgen/$entry
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_word_addrgen/$exit
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_word_addrgen/root_register_req
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_word_addrgen/root_register_ack
      -- 
    ack_1263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_661_final_reg_ack_1, ack => convTranspose_CP_39_elements(151)); -- 
    -- CP-element group 152:  transition  input  output  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	390 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152:  members (6) 
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_664_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_664_Sample/ra
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_664_Update/cr
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_664_Update/$entry
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_664_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_664_update_start_
      -- 
    ra_1272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_664_inst_ack_0, ack => convTranspose_CP_39_elements(152)); -- 
    cr_1276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(152), ack => RPIPE_ConvTranspose_input_pipe_664_inst_req_1); -- 
    -- CP-element group 153:  fork  transition  input  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153: 	156 
    -- CP-element group 153:  members (9) 
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_668_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_664_Update/ca
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_664_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_668_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_664_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_677_Sample/rr
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_677_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_677_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_668_Sample/rr
      -- 
    ca_1277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_664_inst_ack_1, ack => convTranspose_CP_39_elements(153)); -- 
    rr_1285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(153), ack => type_cast_668_inst_req_0); -- 
    rr_1299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(153), ack => RPIPE_ConvTranspose_input_pipe_677_inst_req_0); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_668_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_668_Sample/ra
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_668_Sample/$exit
      -- 
    ra_1286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_668_inst_ack_0, ack => convTranspose_CP_39_elements(154)); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	390 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	184 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_668_Update/ca
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_668_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_668_update_completed_
      -- 
    ca_1291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_668_inst_ack_1, ack => convTranspose_CP_39_elements(155)); -- 
    -- CP-element group 156:  transition  input  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	153 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	157 
    -- CP-element group 156:  members (6) 
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_677_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_677_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_677_Sample/ra
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_677_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_677_update_start_
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_677_sample_completed_
      -- 
    ra_1300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_677_inst_ack_0, ack => convTranspose_CP_39_elements(156)); -- 
    cr_1304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(156), ack => RPIPE_ConvTranspose_input_pipe_677_inst_req_1); -- 
    -- CP-element group 157:  fork  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	156 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157: 	160 
    -- CP-element group 157:  members (9) 
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_695_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_681_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_681_Sample/rr
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_681_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_677_Update/ca
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_677_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_677_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_695_Sample/rr
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_695_Sample/$entry
      -- 
    ca_1305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_677_inst_ack_1, ack => convTranspose_CP_39_elements(157)); -- 
    rr_1313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(157), ack => type_cast_681_inst_req_0); -- 
    rr_1327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(157), ack => RPIPE_ConvTranspose_input_pipe_695_inst_req_0); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_681_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_681_Sample/ra
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_681_Sample/$exit
      -- 
    ra_1314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_681_inst_ack_0, ack => convTranspose_CP_39_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	390 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	184 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_681_Update/ca
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_681_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_681_update_completed_
      -- 
    ca_1319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_681_inst_ack_1, ack => convTranspose_CP_39_elements(159)); -- 
    -- CP-element group 160:  transition  input  output  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	157 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (6) 
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_695_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_695_Update/cr
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_695_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_695_Sample/ra
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_695_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_695_update_start_
      -- 
    ra_1328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_695_inst_ack_0, ack => convTranspose_CP_39_elements(160)); -- 
    cr_1332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(160), ack => RPIPE_ConvTranspose_input_pipe_695_inst_req_1); -- 
    -- CP-element group 161:  fork  transition  input  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161: 	164 
    -- CP-element group 161:  members (9) 
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_713_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_695_Update/ca
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_713_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_695_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_699_Sample/rr
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_699_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_713_Sample/rr
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_695_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_699_sample_start_
      -- 
    ca_1333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_695_inst_ack_1, ack => convTranspose_CP_39_elements(161)); -- 
    rr_1341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(161), ack => type_cast_699_inst_req_0); -- 
    rr_1355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(161), ack => RPIPE_ConvTranspose_input_pipe_713_inst_req_0); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_699_Sample/ra
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_699_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_699_sample_completed_
      -- 
    ra_1342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_699_inst_ack_0, ack => convTranspose_CP_39_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	390 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	184 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_699_Update/ca
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_699_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_699_update_completed_
      -- 
    ca_1347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_699_inst_ack_1, ack => convTranspose_CP_39_elements(163)); -- 
    -- CP-element group 164:  transition  input  output  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	161 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (6) 
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_713_update_start_
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_713_Update/cr
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_713_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_713_Sample/ra
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_713_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_713_sample_completed_
      -- 
    ra_1356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_713_inst_ack_0, ack => convTranspose_CP_39_elements(164)); -- 
    cr_1360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(164), ack => RPIPE_ConvTranspose_input_pipe_713_inst_req_1); -- 
    -- CP-element group 165:  fork  transition  input  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165: 	168 
    -- CP-element group 165:  members (9) 
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_713_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_717_Sample/rr
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_717_Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_717_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_713_Update/ca
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_731_Sample/rr
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_731_Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_713_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_731_sample_start_
      -- 
    ca_1361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_713_inst_ack_1, ack => convTranspose_CP_39_elements(165)); -- 
    rr_1369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(165), ack => type_cast_717_inst_req_0); -- 
    rr_1383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(165), ack => RPIPE_ConvTranspose_input_pipe_731_inst_req_0); -- 
    -- CP-element group 166:  transition  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_717_sample_completed_
      -- CP-element group 166: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_717_Sample/ra
      -- CP-element group 166: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_717_Sample/$exit
      -- 
    ra_1370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_717_inst_ack_0, ack => convTranspose_CP_39_elements(166)); -- 
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	390 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	184 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_717_Update/$exit
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_717_Update/ca
      -- CP-element group 167: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_717_update_completed_
      -- 
    ca_1375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_717_inst_ack_1, ack => convTranspose_CP_39_elements(167)); -- 
    -- CP-element group 168:  transition  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	165 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (6) 
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_731_Update/cr
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_731_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_731_Sample/ra
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_731_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_731_update_start_
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_731_sample_completed_
      -- 
    ra_1384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_731_inst_ack_0, ack => convTranspose_CP_39_elements(168)); -- 
    cr_1388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(168), ack => RPIPE_ConvTranspose_input_pipe_731_inst_req_1); -- 
    -- CP-element group 169:  fork  transition  input  output  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169: 	172 
    -- CP-element group 169:  members (9) 
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_735_Sample/rr
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_749_Sample/$entry
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_749_Sample/rr
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_749_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_735_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_731_Update/ca
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_731_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_731_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_735_Sample/$entry
      -- 
    ca_1389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_731_inst_ack_1, ack => convTranspose_CP_39_elements(169)); -- 
    rr_1397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(169), ack => type_cast_735_inst_req_0); -- 
    rr_1411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(169), ack => RPIPE_ConvTranspose_input_pipe_749_inst_req_0); -- 
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_735_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_735_Sample/ra
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_735_sample_completed_
      -- 
    ra_1398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_735_inst_ack_0, ack => convTranspose_CP_39_elements(170)); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	390 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	184 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_735_Update/ca
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_735_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_735_update_completed_
      -- 
    ca_1403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_735_inst_ack_1, ack => convTranspose_CP_39_elements(171)); -- 
    -- CP-element group 172:  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	169 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (6) 
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_749_Sample/ra
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_749_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_749_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_749_update_start_
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_749_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_749_Update/cr
      -- 
    ra_1412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_749_inst_ack_0, ack => convTranspose_CP_39_elements(172)); -- 
    cr_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(172), ack => RPIPE_ConvTranspose_input_pipe_749_inst_req_1); -- 
    -- CP-element group 173:  fork  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173: 	176 
    -- CP-element group 173:  members (9) 
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_749_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_749_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_749_Update/ca
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_753_sample_start_
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_753_Sample/$entry
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_753_Sample/rr
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_767_sample_start_
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_767_Sample/$entry
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_767_Sample/rr
      -- 
    ca_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_749_inst_ack_1, ack => convTranspose_CP_39_elements(173)); -- 
    rr_1425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(173), ack => type_cast_753_inst_req_0); -- 
    rr_1439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(173), ack => RPIPE_ConvTranspose_input_pipe_767_inst_req_0); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_753_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_753_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_753_Sample/ra
      -- 
    ra_1426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_753_inst_ack_0, ack => convTranspose_CP_39_elements(174)); -- 
    -- CP-element group 175:  transition  input  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	390 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	184 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_753_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_753_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_753_Update/ca
      -- 
    ca_1431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_753_inst_ack_1, ack => convTranspose_CP_39_elements(175)); -- 
    -- CP-element group 176:  transition  input  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	173 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176:  members (6) 
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_767_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_767_update_start_
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_767_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_767_Sample/ra
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_767_Update/$entry
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_767_Update/cr
      -- 
    ra_1440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_767_inst_ack_0, ack => convTranspose_CP_39_elements(176)); -- 
    cr_1444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(176), ack => RPIPE_ConvTranspose_input_pipe_767_inst_req_1); -- 
    -- CP-element group 177:  fork  transition  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177: 	180 
    -- CP-element group 177:  members (9) 
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_767_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_767_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_767_Update/ca
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_771_sample_start_
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_771_Sample/$entry
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_771_Sample/rr
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_785_sample_start_
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_785_Sample/$entry
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_785_Sample/rr
      -- 
    ca_1445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_767_inst_ack_1, ack => convTranspose_CP_39_elements(177)); -- 
    rr_1453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(177), ack => type_cast_771_inst_req_0); -- 
    rr_1467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(177), ack => RPIPE_ConvTranspose_input_pipe_785_inst_req_0); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_771_sample_completed_
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_771_Sample/$exit
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_771_Sample/ra
      -- 
    ra_1454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_771_inst_ack_0, ack => convTranspose_CP_39_elements(178)); -- 
    -- CP-element group 179:  transition  input  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	390 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	184 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_771_update_completed_
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_771_Update/$exit
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_771_Update/ca
      -- 
    ca_1459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_771_inst_ack_1, ack => convTranspose_CP_39_elements(179)); -- 
    -- CP-element group 180:  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	177 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180:  members (6) 
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_785_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_785_update_start_
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_785_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_785_Sample/ra
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_785_Update/$entry
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_785_Update/cr
      -- 
    ra_1468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_785_inst_ack_0, ack => convTranspose_CP_39_elements(180)); -- 
    cr_1472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(180), ack => RPIPE_ConvTranspose_input_pipe_785_inst_req_1); -- 
    -- CP-element group 181:  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (6) 
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_785_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_785_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_785_Update/ca
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_789_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_789_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_789_Sample/rr
      -- 
    ca_1473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_785_inst_ack_1, ack => convTranspose_CP_39_elements(181)); -- 
    rr_1481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(181), ack => type_cast_789_inst_req_0); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_789_sample_completed_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_789_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_789_Sample/ra
      -- 
    ra_1482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_789_inst_ack_0, ack => convTranspose_CP_39_elements(182)); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	390 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_789_update_completed_
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_789_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_789_Update/ca
      -- 
    ca_1487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_789_inst_ack_1, ack => convTranspose_CP_39_elements(183)); -- 
    -- CP-element group 184:  join  transition  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	151 
    -- CP-element group 184: 	155 
    -- CP-element group 184: 	159 
    -- CP-element group 184: 	163 
    -- CP-element group 184: 	167 
    -- CP-element group 184: 	171 
    -- CP-element group 184: 	175 
    -- CP-element group 184: 	179 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (9) 
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Sample/ptr_deref_797_Split/$entry
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Sample/ptr_deref_797_Split/$exit
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Sample/ptr_deref_797_Split/split_req
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Sample/ptr_deref_797_Split/split_ack
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Sample/word_access_start/$entry
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Sample/word_access_start/word_0/$entry
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Sample/word_access_start/word_0/rr
      -- 
    rr_1525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(184), ack => ptr_deref_797_store_0_req_0); -- 
    convTranspose_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(151) & convTranspose_CP_39_elements(155) & convTranspose_CP_39_elements(159) & convTranspose_CP_39_elements(163) & convTranspose_CP_39_elements(167) & convTranspose_CP_39_elements(171) & convTranspose_CP_39_elements(175) & convTranspose_CP_39_elements(179) & convTranspose_CP_39_elements(183);
      gj_convTranspose_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (5) 
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Sample/word_access_start/$exit
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Sample/word_access_start/word_0/$exit
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Sample/word_access_start/word_0/ra
      -- 
    ra_1526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_797_store_0_ack_0, ack => convTranspose_CP_39_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	390 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (5) 
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Update/word_access_complete/$exit
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Update/word_access_complete/word_0/$exit
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Update/word_access_complete/word_0/ca
      -- 
    ca_1537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_797_store_0_ack_1, ack => convTranspose_CP_39_elements(186)); -- 
    -- CP-element group 187:  branch  join  transition  place  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	148 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: 	189 
    -- CP-element group 187:  members (10) 
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810__exit__
      -- CP-element group 187: 	 branch_block_stmt_32/if_stmt_811__entry__
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/$exit
      -- CP-element group 187: 	 branch_block_stmt_32/if_stmt_811_dead_link/$entry
      -- CP-element group 187: 	 branch_block_stmt_32/if_stmt_811_eval_test/$entry
      -- CP-element group 187: 	 branch_block_stmt_32/if_stmt_811_eval_test/$exit
      -- CP-element group 187: 	 branch_block_stmt_32/if_stmt_811_eval_test/branch_req
      -- CP-element group 187: 	 branch_block_stmt_32/R_exitcond2_812_place
      -- CP-element group 187: 	 branch_block_stmt_32/if_stmt_811_if_link/$entry
      -- CP-element group 187: 	 branch_block_stmt_32/if_stmt_811_else_link/$entry
      -- 
    branch_req_1545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(187), ack => if_stmt_811_branch_req_0); -- 
    convTranspose_cp_element_group_187: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_187"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(148) & convTranspose_CP_39_elements(186);
      gj_convTranspose_cp_element_group_187 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(187), clk => clk, reset => reset); --
    end block;
    -- CP-element group 188:  merge  transition  place  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	391 
    -- CP-element group 188:  members (13) 
      -- CP-element group 188: 	 branch_block_stmt_32/merge_stmt_817__exit__
      -- CP-element group 188: 	 branch_block_stmt_32/forx_xend250x_xloopexit_forx_xend250
      -- CP-element group 188: 	 branch_block_stmt_32/merge_stmt_817_PhiAck/dummy
      -- CP-element group 188: 	 branch_block_stmt_32/merge_stmt_817_PhiReqMerge
      -- CP-element group 188: 	 branch_block_stmt_32/forx_xend250x_xloopexit_forx_xend250_PhiReq/$entry
      -- CP-element group 188: 	 branch_block_stmt_32/merge_stmt_817_PhiAck/$entry
      -- CP-element group 188: 	 branch_block_stmt_32/forx_xend250x_xloopexit_forx_xend250_PhiReq/$exit
      -- CP-element group 188: 	 branch_block_stmt_32/if_stmt_811_if_link/$exit
      -- CP-element group 188: 	 branch_block_stmt_32/if_stmt_811_if_link/if_choice_transition
      -- CP-element group 188: 	 branch_block_stmt_32/forx_xbody196_forx_xend250x_xloopexit
      -- CP-element group 188: 	 branch_block_stmt_32/merge_stmt_817_PhiAck/$exit
      -- CP-element group 188: 	 branch_block_stmt_32/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$exit
      -- CP-element group 188: 	 branch_block_stmt_32/forx_xbody196_forx_xend250x_xloopexit_PhiReq/$entry
      -- 
    if_choice_transition_1550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_811_branch_ack_1, ack => convTranspose_CP_39_elements(188)); -- 
    -- CP-element group 189:  fork  transition  place  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	187 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	386 
    -- CP-element group 189: 	387 
    -- CP-element group 189:  members (12) 
      -- CP-element group 189: 	 branch_block_stmt_32/if_stmt_811_else_link/$exit
      -- CP-element group 189: 	 branch_block_stmt_32/if_stmt_811_else_link/else_choice_transition
      -- CP-element group 189: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196
      -- CP-element group 189: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_sources/type_cast_651/SplitProtocol/Update/cr
      -- CP-element group 189: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_sources/type_cast_651/SplitProtocol/Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_sources/type_cast_651/SplitProtocol/Sample/rr
      -- CP-element group 189: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_sources/type_cast_651/SplitProtocol/Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_sources/type_cast_651/SplitProtocol/$entry
      -- CP-element group 189: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_sources/type_cast_651/$entry
      -- CP-element group 189: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_sources/$entry
      -- CP-element group 189: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_648/$entry
      -- CP-element group 189: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/$entry
      -- 
    else_choice_transition_1554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_811_branch_ack_0, ack => convTranspose_CP_39_elements(189)); -- 
    cr_3075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(189), ack => type_cast_651_inst_req_1); -- 
    rr_3070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(189), ack => type_cast_651_inst_req_0); -- 
    -- CP-element group 190:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	391 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190: 	193 
    -- CP-element group 190:  members (18) 
      -- CP-element group 190: 	 branch_block_stmt_32/merge_stmt_842__exit__
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_848_to_assign_stmt_877__entry__
      -- CP-element group 190: 	 branch_block_stmt_32/merge_stmt_842_PhiReqMerge
      -- CP-element group 190: 	 branch_block_stmt_32/if_stmt_836_if_link/$exit
      -- CP-element group 190: 	 branch_block_stmt_32/if_stmt_836_if_link/if_choice_transition
      -- CP-element group 190: 	 branch_block_stmt_32/forx_xend250_bbx_xnph481
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_848_to_assign_stmt_877/$entry
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_848_to_assign_stmt_877/type_cast_863_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_848_to_assign_stmt_877/type_cast_863_update_start_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_848_to_assign_stmt_877/type_cast_863_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_848_to_assign_stmt_877/type_cast_863_Sample/rr
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_848_to_assign_stmt_877/type_cast_863_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_848_to_assign_stmt_877/type_cast_863_Update/cr
      -- CP-element group 190: 	 branch_block_stmt_32/forx_xend250_bbx_xnph481_PhiReq/$entry
      -- CP-element group 190: 	 branch_block_stmt_32/forx_xend250_bbx_xnph481_PhiReq/$exit
      -- CP-element group 190: 	 branch_block_stmt_32/merge_stmt_842_PhiAck/$entry
      -- CP-element group 190: 	 branch_block_stmt_32/merge_stmt_842_PhiAck/$exit
      -- CP-element group 190: 	 branch_block_stmt_32/merge_stmt_842_PhiAck/dummy
      -- 
    if_choice_transition_1572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_836_branch_ack_1, ack => convTranspose_CP_39_elements(190)); -- 
    rr_1589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => type_cast_863_inst_req_0); -- 
    cr_1594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(190), ack => type_cast_863_inst_req_1); -- 
    -- CP-element group 191:  transition  place  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	391 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	398 
    -- CP-element group 191:  members (5) 
      -- CP-element group 191: 	 branch_block_stmt_32/if_stmt_836_else_link/$exit
      -- CP-element group 191: 	 branch_block_stmt_32/if_stmt_836_else_link/else_choice_transition
      -- CP-element group 191: 	 branch_block_stmt_32/forx_xend250_forx_xend273
      -- CP-element group 191: 	 branch_block_stmt_32/forx_xend250_forx_xend273_PhiReq/$exit
      -- CP-element group 191: 	 branch_block_stmt_32/forx_xend250_forx_xend273_PhiReq/$entry
      -- 
    else_choice_transition_1576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_836_branch_ack_0, ack => convTranspose_CP_39_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_848_to_assign_stmt_877/type_cast_863_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_848_to_assign_stmt_877/type_cast_863_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_848_to_assign_stmt_877/type_cast_863_Sample/ra
      -- 
    ra_1590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_863_inst_ack_0, ack => convTranspose_CP_39_elements(192)); -- 
    -- CP-element group 193:  transition  place  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	190 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	392 
    -- CP-element group 193:  members (9) 
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_848_to_assign_stmt_877__exit__
      -- CP-element group 193: 	 branch_block_stmt_32/bbx_xnph481_forx_xbody266
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_848_to_assign_stmt_877/$exit
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_848_to_assign_stmt_877/type_cast_863_update_completed_
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_848_to_assign_stmt_877/type_cast_863_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_848_to_assign_stmt_877/type_cast_863_Update/ca
      -- CP-element group 193: 	 branch_block_stmt_32/bbx_xnph481_forx_xbody266_PhiReq/$entry
      -- CP-element group 193: 	 branch_block_stmt_32/bbx_xnph481_forx_xbody266_PhiReq/phi_stmt_880/$entry
      -- CP-element group 193: 	 branch_block_stmt_32/bbx_xnph481_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_sources/$entry
      -- 
    ca_1595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_863_inst_ack_1, ack => convTranspose_CP_39_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	397 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	200 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_final_index_sum_regn_sample_complete
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_final_index_sum_regn_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_final_index_sum_regn_Sample/ack
      -- 
    ack_1624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_892_index_offset_ack_0, ack => convTranspose_CP_39_elements(194)); -- 
    -- CP-element group 195:  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	397 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (11) 
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/addr_of_893_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_root_address_calculated
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_offset_calculated
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_final_index_sum_regn_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_final_index_sum_regn_Update/ack
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_base_plus_offset/$entry
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_base_plus_offset/$exit
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_base_plus_offset/sum_rename_req
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_base_plus_offset/sum_rename_ack
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/addr_of_893_request/$entry
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/addr_of_893_request/req
      -- 
    ack_1629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_892_index_offset_ack_1, ack => convTranspose_CP_39_elements(195)); -- 
    req_1638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(195), ack => addr_of_893_final_reg_req_0); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/addr_of_893_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/addr_of_893_request/$exit
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/addr_of_893_request/ack
      -- 
    ack_1639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_893_final_reg_ack_0, ack => convTranspose_CP_39_elements(196)); -- 
    -- CP-element group 197:  join  fork  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	397 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (28) 
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/addr_of_893_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/addr_of_893_complete/$exit
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/addr_of_893_complete/ack
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_sample_start_
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_base_address_calculated
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_word_address_calculated
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_root_address_calculated
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_base_address_resized
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_base_addr_resize/$entry
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_base_addr_resize/$exit
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_base_addr_resize/base_resize_req
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_base_addr_resize/base_resize_ack
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_base_plus_offset/$entry
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_base_plus_offset/$exit
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_base_plus_offset/sum_rename_req
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_base_plus_offset/sum_rename_ack
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_word_addrgen/$entry
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_word_addrgen/$exit
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_word_addrgen/root_register_req
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_word_addrgen/root_register_ack
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Sample/$entry
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Sample/ptr_deref_896_Split/$entry
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Sample/ptr_deref_896_Split/$exit
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Sample/ptr_deref_896_Split/split_req
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Sample/ptr_deref_896_Split/split_ack
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Sample/word_access_start/$entry
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Sample/word_access_start/word_0/$entry
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Sample/word_access_start/word_0/rr
      -- 
    ack_1644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_893_final_reg_ack_1, ack => convTranspose_CP_39_elements(197)); -- 
    rr_1682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(197), ack => ptr_deref_896_store_0_req_0); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198:  members (5) 
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Sample/word_access_start/$exit
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Sample/word_access_start/word_0/$exit
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Sample/word_access_start/word_0/ra
      -- 
    ra_1683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_896_store_0_ack_0, ack => convTranspose_CP_39_elements(198)); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	397 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (5) 
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Update/word_access_complete/$exit
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Update/word_access_complete/word_0/$exit
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Update/word_access_complete/word_0/ca
      -- 
    ca_1694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_896_store_0_ack_1, ack => convTranspose_CP_39_elements(199)); -- 
    -- CP-element group 200:  branch  join  transition  place  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	194 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200: 	202 
    -- CP-element group 200:  members (10) 
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910__exit__
      -- CP-element group 200: 	 branch_block_stmt_32/if_stmt_911__entry__
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/$exit
      -- CP-element group 200: 	 branch_block_stmt_32/if_stmt_911_dead_link/$entry
      -- CP-element group 200: 	 branch_block_stmt_32/if_stmt_911_eval_test/$entry
      -- CP-element group 200: 	 branch_block_stmt_32/if_stmt_911_eval_test/$exit
      -- CP-element group 200: 	 branch_block_stmt_32/if_stmt_911_eval_test/branch_req
      -- CP-element group 200: 	 branch_block_stmt_32/R_exitcond_912_place
      -- CP-element group 200: 	 branch_block_stmt_32/if_stmt_911_if_link/$entry
      -- CP-element group 200: 	 branch_block_stmt_32/if_stmt_911_else_link/$entry
      -- 
    branch_req_1702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(200), ack => if_stmt_911_branch_req_0); -- 
    convTranspose_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(194) & convTranspose_CP_39_elements(199);
      gj_convTranspose_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  merge  transition  place  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	398 
    -- CP-element group 201:  members (13) 
      -- CP-element group 201: 	 branch_block_stmt_32/merge_stmt_917__exit__
      -- CP-element group 201: 	 branch_block_stmt_32/forx_xend273x_xloopexit_forx_xend273
      -- CP-element group 201: 	 branch_block_stmt_32/merge_stmt_917_PhiReqMerge
      -- CP-element group 201: 	 branch_block_stmt_32/if_stmt_911_if_link/$exit
      -- CP-element group 201: 	 branch_block_stmt_32/if_stmt_911_if_link/if_choice_transition
      -- CP-element group 201: 	 branch_block_stmt_32/forx_xbody266_forx_xend273x_xloopexit
      -- CP-element group 201: 	 branch_block_stmt_32/forx_xend273x_xloopexit_forx_xend273_PhiReq/$exit
      -- CP-element group 201: 	 branch_block_stmt_32/forx_xend273x_xloopexit_forx_xend273_PhiReq/$entry
      -- CP-element group 201: 	 branch_block_stmt_32/merge_stmt_917_PhiAck/dummy
      -- CP-element group 201: 	 branch_block_stmt_32/merge_stmt_917_PhiAck/$exit
      -- CP-element group 201: 	 branch_block_stmt_32/merge_stmt_917_PhiAck/$entry
      -- CP-element group 201: 	 branch_block_stmt_32/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$exit
      -- CP-element group 201: 	 branch_block_stmt_32/forx_xbody266_forx_xend273x_xloopexit_PhiReq/$entry
      -- 
    if_choice_transition_1707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_911_branch_ack_1, ack => convTranspose_CP_39_elements(201)); -- 
    -- CP-element group 202:  fork  transition  place  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	200 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	393 
    -- CP-element group 202: 	394 
    -- CP-element group 202:  members (12) 
      -- CP-element group 202: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_sources/type_cast_883/SplitProtocol/Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_32/if_stmt_911_else_link/$exit
      -- CP-element group 202: 	 branch_block_stmt_32/if_stmt_911_else_link/else_choice_transition
      -- CP-element group 202: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266
      -- CP-element group 202: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_sources/type_cast_883/SplitProtocol/$entry
      -- CP-element group 202: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_sources/type_cast_883/$entry
      -- CP-element group 202: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_sources/$entry
      -- CP-element group 202: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_880/$entry
      -- CP-element group 202: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/$entry
      -- CP-element group 202: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_sources/type_cast_883/SplitProtocol/Update/cr
      -- CP-element group 202: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_sources/type_cast_883/SplitProtocol/Update/$entry
      -- CP-element group 202: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_sources/type_cast_883/SplitProtocol/Sample/rr
      -- 
    else_choice_transition_1711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_911_branch_ack_0, ack => convTranspose_CP_39_elements(202)); -- 
    cr_3152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(202), ack => type_cast_883_inst_req_1); -- 
    rr_3147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(202), ack => type_cast_883_inst_req_0); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	398 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/call_stmt_922_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/call_stmt_922_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/call_stmt_922_Sample/cra
      -- 
    cra_1725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_922_call_ack_0, ack => convTranspose_CP_39_elements(203)); -- 
    -- CP-element group 204:  transition  input  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	398 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (6) 
      -- CP-element group 204: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/call_stmt_922_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/call_stmt_922_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/call_stmt_922_Update/cca
      -- CP-element group 204: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/type_cast_927_sample_start_
      -- CP-element group 204: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/type_cast_927_Sample/$entry
      -- CP-element group 204: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/type_cast_927_Sample/rr
      -- 
    cca_1730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_922_call_ack_1, ack => convTranspose_CP_39_elements(204)); -- 
    rr_1738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(204), ack => type_cast_927_inst_req_0); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/type_cast_927_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/type_cast_927_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/type_cast_927_Sample/ra
      -- 
    ra_1739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_927_inst_ack_0, ack => convTranspose_CP_39_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	398 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	319 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/type_cast_927_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/type_cast_927_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/type_cast_927_Update/ca
      -- 
    ca_1744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_927_inst_ack_1, ack => convTranspose_CP_39_elements(206)); -- 
    -- CP-element group 207:  transition  input  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	398 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (6) 
      -- CP-element group 207: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_929_sample_completed_
      -- CP-element group 207: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_929_update_start_
      -- CP-element group 207: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_929_Sample/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_929_Sample/ack
      -- CP-element group 207: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_929_Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_929_Update/req
      -- 
    ack_1753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_929_inst_ack_0, ack => convTranspose_CP_39_elements(207)); -- 
    req_1757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(207), ack => WPIPE_Block0_start_929_inst_req_1); -- 
    -- CP-element group 208:  transition  input  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208:  members (6) 
      -- CP-element group 208: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_929_update_completed_
      -- CP-element group 208: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_929_Update/$exit
      -- CP-element group 208: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_929_Update/ack
      -- CP-element group 208: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_932_sample_start_
      -- CP-element group 208: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_932_Sample/$entry
      -- CP-element group 208: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_932_Sample/req
      -- 
    ack_1758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_929_inst_ack_1, ack => convTranspose_CP_39_elements(208)); -- 
    req_1766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(208), ack => WPIPE_Block0_start_932_inst_req_0); -- 
    -- CP-element group 209:  transition  input  output  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209:  members (6) 
      -- CP-element group 209: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_932_sample_completed_
      -- CP-element group 209: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_932_update_start_
      -- CP-element group 209: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_932_Sample/$exit
      -- CP-element group 209: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_932_Sample/ack
      -- CP-element group 209: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_932_Update/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_932_Update/req
      -- 
    ack_1767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_932_inst_ack_0, ack => convTranspose_CP_39_elements(209)); -- 
    req_1771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(209), ack => WPIPE_Block0_start_932_inst_req_1); -- 
    -- CP-element group 210:  transition  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210:  members (6) 
      -- CP-element group 210: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_932_update_completed_
      -- CP-element group 210: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_932_Update/$exit
      -- CP-element group 210: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_932_Update/ack
      -- CP-element group 210: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_935_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_935_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_935_Sample/req
      -- 
    ack_1772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_932_inst_ack_1, ack => convTranspose_CP_39_elements(210)); -- 
    req_1780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(210), ack => WPIPE_Block0_start_935_inst_req_0); -- 
    -- CP-element group 211:  transition  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	212 
    -- CP-element group 211:  members (6) 
      -- CP-element group 211: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_935_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_935_update_start_
      -- CP-element group 211: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_935_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_935_Sample/ack
      -- CP-element group 211: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_935_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_935_Update/req
      -- 
    ack_1781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_935_inst_ack_0, ack => convTranspose_CP_39_elements(211)); -- 
    req_1785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(211), ack => WPIPE_Block0_start_935_inst_req_1); -- 
    -- CP-element group 212:  transition  input  output  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	211 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	213 
    -- CP-element group 212:  members (6) 
      -- CP-element group 212: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_935_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_935_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_935_Update/ack
      -- CP-element group 212: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_938_sample_start_
      -- CP-element group 212: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_938_Sample/$entry
      -- CP-element group 212: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_938_Sample/req
      -- 
    ack_1786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_935_inst_ack_1, ack => convTranspose_CP_39_elements(212)); -- 
    req_1794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(212), ack => WPIPE_Block0_start_938_inst_req_0); -- 
    -- CP-element group 213:  transition  input  output  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	212 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213:  members (6) 
      -- CP-element group 213: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_938_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_938_update_start_
      -- CP-element group 213: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_938_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_938_Sample/ack
      -- CP-element group 213: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_938_Update/$entry
      -- CP-element group 213: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_938_Update/req
      -- 
    ack_1795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_938_inst_ack_0, ack => convTranspose_CP_39_elements(213)); -- 
    req_1799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(213), ack => WPIPE_Block0_start_938_inst_req_1); -- 
    -- CP-element group 214:  transition  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	213 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (6) 
      -- CP-element group 214: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_938_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_938_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_938_Update/ack
      -- CP-element group 214: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_941_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_941_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_941_Sample/req
      -- 
    ack_1800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_938_inst_ack_1, ack => convTranspose_CP_39_elements(214)); -- 
    req_1808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(214), ack => WPIPE_Block0_start_941_inst_req_0); -- 
    -- CP-element group 215:  transition  input  output  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215:  members (6) 
      -- CP-element group 215: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_941_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_941_update_start_
      -- CP-element group 215: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_941_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_941_Sample/ack
      -- CP-element group 215: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_941_Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_941_Update/req
      -- 
    ack_1809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_941_inst_ack_0, ack => convTranspose_CP_39_elements(215)); -- 
    req_1813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(215), ack => WPIPE_Block0_start_941_inst_req_1); -- 
    -- CP-element group 216:  transition  input  output  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (6) 
      -- CP-element group 216: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_941_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_941_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_941_Update/ack
      -- CP-element group 216: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_944_sample_start_
      -- CP-element group 216: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_944_Sample/$entry
      -- CP-element group 216: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_944_Sample/req
      -- 
    ack_1814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_941_inst_ack_1, ack => convTranspose_CP_39_elements(216)); -- 
    req_1822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(216), ack => WPIPE_Block0_start_944_inst_req_0); -- 
    -- CP-element group 217:  transition  input  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (6) 
      -- CP-element group 217: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_944_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_944_update_start_
      -- CP-element group 217: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_944_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_944_Sample/ack
      -- CP-element group 217: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_944_Update/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_944_Update/req
      -- 
    ack_1823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_944_inst_ack_0, ack => convTranspose_CP_39_elements(217)); -- 
    req_1827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(217), ack => WPIPE_Block0_start_944_inst_req_1); -- 
    -- CP-element group 218:  transition  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (6) 
      -- CP-element group 218: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_944_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_944_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_944_Update/ack
      -- CP-element group 218: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_947_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_947_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_947_Sample/req
      -- 
    ack_1828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_944_inst_ack_1, ack => convTranspose_CP_39_elements(218)); -- 
    req_1836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(218), ack => WPIPE_Block0_start_947_inst_req_0); -- 
    -- CP-element group 219:  transition  input  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219:  members (6) 
      -- CP-element group 219: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_947_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_947_update_start_
      -- CP-element group 219: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_947_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_947_Sample/ack
      -- CP-element group 219: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_947_Update/$entry
      -- CP-element group 219: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_947_Update/req
      -- 
    ack_1837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_947_inst_ack_0, ack => convTranspose_CP_39_elements(219)); -- 
    req_1841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(219), ack => WPIPE_Block0_start_947_inst_req_1); -- 
    -- CP-element group 220:  transition  input  output  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	221 
    -- CP-element group 220:  members (6) 
      -- CP-element group 220: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_947_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_947_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_947_Update/ack
      -- CP-element group 220: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_950_sample_start_
      -- CP-element group 220: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_950_Sample/$entry
      -- CP-element group 220: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_950_Sample/req
      -- 
    ack_1842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_947_inst_ack_1, ack => convTranspose_CP_39_elements(220)); -- 
    req_1850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(220), ack => WPIPE_Block0_start_950_inst_req_0); -- 
    -- CP-element group 221:  transition  input  output  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	220 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	222 
    -- CP-element group 221:  members (6) 
      -- CP-element group 221: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_950_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_950_update_start_
      -- CP-element group 221: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_950_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_950_Sample/ack
      -- CP-element group 221: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_950_Update/$entry
      -- CP-element group 221: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_950_Update/req
      -- 
    ack_1851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_950_inst_ack_0, ack => convTranspose_CP_39_elements(221)); -- 
    req_1855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(221), ack => WPIPE_Block0_start_950_inst_req_1); -- 
    -- CP-element group 222:  transition  input  output  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	221 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (6) 
      -- CP-element group 222: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_950_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_950_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_950_Update/ack
      -- CP-element group 222: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_953_sample_start_
      -- CP-element group 222: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_953_Sample/$entry
      -- CP-element group 222: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_953_Sample/req
      -- 
    ack_1856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_950_inst_ack_1, ack => convTranspose_CP_39_elements(222)); -- 
    req_1864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(222), ack => WPIPE_Block0_start_953_inst_req_0); -- 
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (6) 
      -- CP-element group 223: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_953_sample_completed_
      -- CP-element group 223: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_953_update_start_
      -- CP-element group 223: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_953_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_953_Sample/ack
      -- CP-element group 223: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_953_Update/$entry
      -- CP-element group 223: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_953_Update/req
      -- 
    ack_1865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_953_inst_ack_0, ack => convTranspose_CP_39_elements(223)); -- 
    req_1869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(223), ack => WPIPE_Block0_start_953_inst_req_1); -- 
    -- CP-element group 224:  transition  input  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	225 
    -- CP-element group 224:  members (6) 
      -- CP-element group 224: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_953_update_completed_
      -- CP-element group 224: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_953_Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_953_Update/ack
      -- CP-element group 224: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_956_sample_start_
      -- CP-element group 224: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_956_Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_956_Sample/req
      -- 
    ack_1870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_953_inst_ack_1, ack => convTranspose_CP_39_elements(224)); -- 
    req_1878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(224), ack => WPIPE_Block0_start_956_inst_req_0); -- 
    -- CP-element group 225:  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	224 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (6) 
      -- CP-element group 225: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_956_sample_completed_
      -- CP-element group 225: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_956_update_start_
      -- CP-element group 225: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_956_Sample/$exit
      -- CP-element group 225: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_956_Sample/ack
      -- CP-element group 225: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_956_Update/$entry
      -- CP-element group 225: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_956_Update/req
      -- 
    ack_1879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_956_inst_ack_0, ack => convTranspose_CP_39_elements(225)); -- 
    req_1883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(225), ack => WPIPE_Block0_start_956_inst_req_1); -- 
    -- CP-element group 226:  transition  input  output  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (6) 
      -- CP-element group 226: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_956_update_completed_
      -- CP-element group 226: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_956_Update/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_956_Update/ack
      -- CP-element group 226: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_960_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_960_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_960_Sample/req
      -- 
    ack_1884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_956_inst_ack_1, ack => convTranspose_CP_39_elements(226)); -- 
    req_1892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(226), ack => WPIPE_Block0_start_960_inst_req_0); -- 
    -- CP-element group 227:  transition  input  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (6) 
      -- CP-element group 227: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_960_sample_completed_
      -- CP-element group 227: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_960_update_start_
      -- CP-element group 227: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_960_Sample/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_960_Sample/ack
      -- CP-element group 227: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_960_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_960_Update/req
      -- 
    ack_1893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_960_inst_ack_0, ack => convTranspose_CP_39_elements(227)); -- 
    req_1897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(227), ack => WPIPE_Block0_start_960_inst_req_1); -- 
    -- CP-element group 228:  transition  input  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228:  members (6) 
      -- CP-element group 228: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_960_update_completed_
      -- CP-element group 228: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_960_Update/$exit
      -- CP-element group 228: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_960_Update/ack
      -- CP-element group 228: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_963_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_963_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_963_Sample/req
      -- 
    ack_1898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_960_inst_ack_1, ack => convTranspose_CP_39_elements(228)); -- 
    req_1906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(228), ack => WPIPE_Block0_start_963_inst_req_0); -- 
    -- CP-element group 229:  transition  input  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (6) 
      -- CP-element group 229: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_963_sample_completed_
      -- CP-element group 229: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_963_update_start_
      -- CP-element group 229: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_963_Sample/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_963_Sample/ack
      -- CP-element group 229: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_963_Update/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_963_Update/req
      -- 
    ack_1907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_963_inst_ack_0, ack => convTranspose_CP_39_elements(229)); -- 
    req_1911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(229), ack => WPIPE_Block0_start_963_inst_req_1); -- 
    -- CP-element group 230:  transition  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (6) 
      -- CP-element group 230: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_963_update_completed_
      -- CP-element group 230: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_963_Update/$exit
      -- CP-element group 230: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_963_Update/ack
      -- CP-element group 230: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_966_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_966_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_966_Sample/req
      -- 
    ack_1912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_963_inst_ack_1, ack => convTranspose_CP_39_elements(230)); -- 
    req_1920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(230), ack => WPIPE_Block0_start_966_inst_req_0); -- 
    -- CP-element group 231:  transition  input  output  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (6) 
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_966_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_966_update_start_
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_966_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_966_Sample/ack
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_966_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_966_Update/req
      -- 
    ack_1921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_966_inst_ack_0, ack => convTranspose_CP_39_elements(231)); -- 
    req_1925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(231), ack => WPIPE_Block0_start_966_inst_req_1); -- 
    -- CP-element group 232:  transition  input  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	319 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_966_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_966_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_966_Update/ack
      -- 
    ack_1926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_966_inst_ack_1, ack => convTranspose_CP_39_elements(232)); -- 
    -- CP-element group 233:  transition  input  output  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	398 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	234 
    -- CP-element group 233:  members (6) 
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_969_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_969_update_start_
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_969_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_969_Sample/ack
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_969_Update/$entry
      -- CP-element group 233: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_969_Update/req
      -- 
    ack_1935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_969_inst_ack_0, ack => convTranspose_CP_39_elements(233)); -- 
    req_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(233), ack => WPIPE_Block1_start_969_inst_req_1); -- 
    -- CP-element group 234:  transition  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	233 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234:  members (6) 
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_969_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_969_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_969_Update/ack
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_972_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_972_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_972_Sample/req
      -- 
    ack_1940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_969_inst_ack_1, ack => convTranspose_CP_39_elements(234)); -- 
    req_1948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(234), ack => WPIPE_Block1_start_972_inst_req_0); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_972_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_972_update_start_
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_972_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_972_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_972_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_972_Update/req
      -- 
    ack_1949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_972_inst_ack_0, ack => convTranspose_CP_39_elements(235)); -- 
    req_1953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(235), ack => WPIPE_Block1_start_972_inst_req_1); -- 
    -- CP-element group 236:  transition  input  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_972_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_972_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_972_Update/ack
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_975_sample_start_
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_975_Sample/$entry
      -- CP-element group 236: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_975_Sample/req
      -- 
    ack_1954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_972_inst_ack_1, ack => convTranspose_CP_39_elements(236)); -- 
    req_1962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(236), ack => WPIPE_Block1_start_975_inst_req_0); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_975_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_975_update_start_
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_975_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_975_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_975_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_975_Update/req
      -- 
    ack_1963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_975_inst_ack_0, ack => convTranspose_CP_39_elements(237)); -- 
    req_1967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(237), ack => WPIPE_Block1_start_975_inst_req_1); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_975_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_975_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_975_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_978_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_978_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_978_Sample/req
      -- 
    ack_1968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_975_inst_ack_1, ack => convTranspose_CP_39_elements(238)); -- 
    req_1976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(238), ack => WPIPE_Block1_start_978_inst_req_0); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_978_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_978_update_start_
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_978_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_978_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_978_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_978_Update/req
      -- 
    ack_1977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_978_inst_ack_0, ack => convTranspose_CP_39_elements(239)); -- 
    req_1981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(239), ack => WPIPE_Block1_start_978_inst_req_1); -- 
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_978_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_978_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_978_Update/ack
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_981_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_981_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_981_Sample/req
      -- 
    ack_1982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_978_inst_ack_1, ack => convTranspose_CP_39_elements(240)); -- 
    req_1990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(240), ack => WPIPE_Block1_start_981_inst_req_0); -- 
    -- CP-element group 241:  transition  input  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_981_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_981_update_start_
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_981_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_981_Sample/ack
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_981_Update/$entry
      -- CP-element group 241: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_981_Update/req
      -- 
    ack_1991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_981_inst_ack_0, ack => convTranspose_CP_39_elements(241)); -- 
    req_1995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(241), ack => WPIPE_Block1_start_981_inst_req_1); -- 
    -- CP-element group 242:  transition  input  output  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (6) 
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_981_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_981_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_981_Update/ack
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_984_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_984_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_984_Sample/req
      -- 
    ack_1996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_981_inst_ack_1, ack => convTranspose_CP_39_elements(242)); -- 
    req_2004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(242), ack => WPIPE_Block1_start_984_inst_req_0); -- 
    -- CP-element group 243:  transition  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (6) 
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_984_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_984_update_start_
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_984_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_984_Sample/ack
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_984_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_984_Update/req
      -- 
    ack_2005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_984_inst_ack_0, ack => convTranspose_CP_39_elements(243)); -- 
    req_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(243), ack => WPIPE_Block1_start_984_inst_req_1); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_987_Sample/req
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_987_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_984_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_984_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_984_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_987_sample_start_
      -- 
    ack_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_984_inst_ack_1, ack => convTranspose_CP_39_elements(244)); -- 
    req_2018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(244), ack => WPIPE_Block1_start_987_inst_req_0); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_987_Update/req
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_987_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_987_Sample/ack
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_987_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_987_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_987_update_start_
      -- 
    ack_2019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_987_inst_ack_0, ack => convTranspose_CP_39_elements(245)); -- 
    req_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(245), ack => WPIPE_Block1_start_987_inst_req_1); -- 
    -- CP-element group 246:  transition  input  output  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (6) 
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_987_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_990_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_990_Sample/req
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_990_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_987_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_987_update_completed_
      -- 
    ack_2024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_987_inst_ack_1, ack => convTranspose_CP_39_elements(246)); -- 
    req_2032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(246), ack => WPIPE_Block1_start_990_inst_req_0); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_990_update_start_
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_990_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_990_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_990_Sample/ack
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_990_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_990_Update/req
      -- 
    ack_2033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_990_inst_ack_0, ack => convTranspose_CP_39_elements(247)); -- 
    req_2037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(247), ack => WPIPE_Block1_start_990_inst_req_1); -- 
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_990_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_990_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_993_Sample/req
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_993_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_993_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_990_Update/ack
      -- 
    ack_2038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_990_inst_ack_1, ack => convTranspose_CP_39_elements(248)); -- 
    req_2046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(248), ack => WPIPE_Block1_start_993_inst_req_0); -- 
    -- CP-element group 249:  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (6) 
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_993_Update/req
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_993_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_993_Sample/ack
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_993_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_993_update_start_
      -- CP-element group 249: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_993_sample_completed_
      -- 
    ack_2047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_993_inst_ack_0, ack => convTranspose_CP_39_elements(249)); -- 
    req_2051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(249), ack => WPIPE_Block1_start_993_inst_req_1); -- 
    -- CP-element group 250:  transition  input  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (6) 
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_996_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_993_Update/ack
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_993_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_996_Sample/req
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_996_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_993_update_completed_
      -- 
    ack_2052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_993_inst_ack_1, ack => convTranspose_CP_39_elements(250)); -- 
    req_2060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(250), ack => WPIPE_Block1_start_996_inst_req_0); -- 
    -- CP-element group 251:  transition  input  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_996_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_996_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_996_update_start_
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_996_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_996_Sample/ack
      -- CP-element group 251: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_996_Update/req
      -- 
    ack_2061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_996_inst_ack_0, ack => convTranspose_CP_39_elements(251)); -- 
    req_2065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(251), ack => WPIPE_Block1_start_996_inst_req_1); -- 
    -- CP-element group 252:  transition  input  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (6) 
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_996_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_999_Sample/req
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_999_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_999_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_996_Update/ack
      -- CP-element group 252: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_996_Update/$exit
      -- 
    ack_2066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_996_inst_ack_1, ack => convTranspose_CP_39_elements(252)); -- 
    req_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(252), ack => WPIPE_Block1_start_999_inst_req_0); -- 
    -- CP-element group 253:  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_999_Update/req
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_999_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_999_Sample/ack
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_999_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_999_update_start_
      -- CP-element group 253: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_999_sample_completed_
      -- 
    ack_2075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_999_inst_ack_0, ack => convTranspose_CP_39_elements(253)); -- 
    req_2079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(253), ack => WPIPE_Block1_start_999_inst_req_1); -- 
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (6) 
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1002_Sample/req
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1002_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1002_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_999_Update/ack
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_999_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_999_update_completed_
      -- 
    ack_2080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_999_inst_ack_1, ack => convTranspose_CP_39_elements(254)); -- 
    req_2088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(254), ack => WPIPE_Block1_start_1002_inst_req_0); -- 
    -- CP-element group 255:  transition  input  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (6) 
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1002_Sample/ack
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1002_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1002_Update/req
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1002_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1002_update_start_
      -- CP-element group 255: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1002_sample_completed_
      -- 
    ack_2089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1002_inst_ack_0, ack => convTranspose_CP_39_elements(255)); -- 
    req_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(255), ack => WPIPE_Block1_start_1002_inst_req_1); -- 
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1002_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1005_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1005_Sample/req
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1002_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1005_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1002_update_completed_
      -- 
    ack_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1002_inst_ack_1, ack => convTranspose_CP_39_elements(256)); -- 
    req_2102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(256), ack => WPIPE_Block1_start_1005_inst_req_0); -- 
    -- CP-element group 257:  transition  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (6) 
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1005_Sample/ack
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1005_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1005_Update/req
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1005_update_start_
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1005_sample_completed_
      -- CP-element group 257: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1005_Sample/$exit
      -- 
    ack_2103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1005_inst_ack_0, ack => convTranspose_CP_39_elements(257)); -- 
    req_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(257), ack => WPIPE_Block1_start_1005_inst_req_1); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	319 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1005_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1005_update_completed_
      -- CP-element group 258: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_1005_Update/ack
      -- 
    ack_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1005_inst_ack_1, ack => convTranspose_CP_39_elements(258)); -- 
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	398 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1008_update_start_
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1008_sample_completed_
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1008_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1008_Update/req
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1008_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1008_Sample/ack
      -- 
    ack_2117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1008_inst_ack_0, ack => convTranspose_CP_39_elements(259)); -- 
    req_2121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(259), ack => WPIPE_Block2_start_1008_inst_req_1); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1011_Sample/req
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1011_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1008_update_completed_
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1011_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1008_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1008_Update/$exit
      -- 
    ack_2122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1008_inst_ack_1, ack => convTranspose_CP_39_elements(260)); -- 
    req_2130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(260), ack => WPIPE_Block2_start_1011_inst_req_0); -- 
    -- CP-element group 261:  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (6) 
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1011_Update/req
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1011_Sample/ack
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1011_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1011_Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1011_update_start_
      -- CP-element group 261: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1011_sample_completed_
      -- 
    ack_2131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1011_inst_ack_0, ack => convTranspose_CP_39_elements(261)); -- 
    req_2135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(261), ack => WPIPE_Block2_start_1011_inst_req_1); -- 
    -- CP-element group 262:  transition  input  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262:  members (6) 
      -- CP-element group 262: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1011_Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1011_update_completed_
      -- CP-element group 262: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1011_Update/ack
      -- CP-element group 262: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1014_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1014_Sample/req
      -- CP-element group 262: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1014_Sample/$entry
      -- 
    ack_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1011_inst_ack_1, ack => convTranspose_CP_39_elements(262)); -- 
    req_2144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(262), ack => WPIPE_Block2_start_1014_inst_req_0); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1014_Update/req
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1014_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1014_Sample/ack
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1014_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1014_update_start_
      -- CP-element group 263: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1014_sample_completed_
      -- 
    ack_2145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1014_inst_ack_0, ack => convTranspose_CP_39_elements(263)); -- 
    req_2149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(263), ack => WPIPE_Block2_start_1014_inst_req_1); -- 
    -- CP-element group 264:  transition  input  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1017_Sample/req
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1017_Sample/$entry
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1017_sample_start_
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1014_Update/ack
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1014_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1014_update_completed_
      -- 
    ack_2150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1014_inst_ack_1, ack => convTranspose_CP_39_elements(264)); -- 
    req_2158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(264), ack => WPIPE_Block2_start_1017_inst_req_0); -- 
    -- CP-element group 265:  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (6) 
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1017_Update/req
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1017_Update/$entry
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1017_Sample/ack
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1017_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1017_update_start_
      -- CP-element group 265: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1017_sample_completed_
      -- 
    ack_2159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1017_inst_ack_0, ack => convTranspose_CP_39_elements(265)); -- 
    req_2163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(265), ack => WPIPE_Block2_start_1017_inst_req_1); -- 
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1020_Sample/req
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1020_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1020_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1017_Update/ack
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1017_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1017_update_completed_
      -- 
    ack_2164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1017_inst_ack_1, ack => convTranspose_CP_39_elements(266)); -- 
    req_2172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(266), ack => WPIPE_Block2_start_1020_inst_req_0); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1020_Update/req
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1020_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1020_Sample/ack
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1020_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1020_update_start_
      -- CP-element group 267: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1020_sample_completed_
      -- 
    ack_2173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1020_inst_ack_0, ack => convTranspose_CP_39_elements(267)); -- 
    req_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(267), ack => WPIPE_Block2_start_1020_inst_req_1); -- 
    -- CP-element group 268:  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (6) 
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1023_Sample/req
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1023_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1023_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1020_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1020_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1020_update_completed_
      -- 
    ack_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1020_inst_ack_1, ack => convTranspose_CP_39_elements(268)); -- 
    req_2186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(268), ack => WPIPE_Block2_start_1023_inst_req_0); -- 
    -- CP-element group 269:  transition  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (6) 
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1023_Update/req
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1023_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1023_Sample/ack
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1023_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1023_update_start_
      -- CP-element group 269: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1023_sample_completed_
      -- 
    ack_2187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1023_inst_ack_0, ack => convTranspose_CP_39_elements(269)); -- 
    req_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(269), ack => WPIPE_Block2_start_1023_inst_req_1); -- 
    -- CP-element group 270:  transition  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1023_Update/ack
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1026_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1026_Sample/req
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1026_Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1023_Update/$exit
      -- CP-element group 270: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1023_update_completed_
      -- 
    ack_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1023_inst_ack_1, ack => convTranspose_CP_39_elements(270)); -- 
    req_2200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(270), ack => WPIPE_Block2_start_1026_inst_req_0); -- 
    -- CP-element group 271:  transition  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (6) 
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1026_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1026_update_start_
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1026_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1026_sample_completed_
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1026_Update/req
      -- CP-element group 271: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1026_Sample/ack
      -- 
    ack_2201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1026_inst_ack_0, ack => convTranspose_CP_39_elements(271)); -- 
    req_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(271), ack => WPIPE_Block2_start_1026_inst_req_1); -- 
    -- CP-element group 272:  transition  input  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (6) 
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1029_Sample/$entry
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1029_Sample/req
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1029_sample_start_
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1026_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1026_update_completed_
      -- CP-element group 272: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1026_Update/ack
      -- 
    ack_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1026_inst_ack_1, ack => convTranspose_CP_39_elements(272)); -- 
    req_2214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(272), ack => WPIPE_Block2_start_1029_inst_req_0); -- 
    -- CP-element group 273:  transition  input  output  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (6) 
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1029_Update/$entry
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1029_Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1029_Sample/ack
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1029_sample_completed_
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1029_update_start_
      -- CP-element group 273: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1029_Update/req
      -- 
    ack_2215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1029_inst_ack_0, ack => convTranspose_CP_39_elements(273)); -- 
    req_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(273), ack => WPIPE_Block2_start_1029_inst_req_1); -- 
    -- CP-element group 274:  transition  input  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (6) 
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1029_update_completed_
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1029_Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1029_Update/ack
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1032_sample_start_
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1032_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1032_Sample/req
      -- 
    ack_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1029_inst_ack_1, ack => convTranspose_CP_39_elements(274)); -- 
    req_2228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(274), ack => WPIPE_Block2_start_1032_inst_req_0); -- 
    -- CP-element group 275:  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1032_sample_completed_
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1032_update_start_
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1032_Update/req
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1032_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1032_Sample/ack
      -- CP-element group 275: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1032_Update/$entry
      -- 
    ack_2229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1032_inst_ack_0, ack => convTranspose_CP_39_elements(275)); -- 
    req_2233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(275), ack => WPIPE_Block2_start_1032_inst_req_1); -- 
    -- CP-element group 276:  transition  input  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (6) 
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1032_update_completed_
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1032_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1035_Sample/req
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1035_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1035_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1032_Update/ack
      -- 
    ack_2234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1032_inst_ack_1, ack => convTranspose_CP_39_elements(276)); -- 
    req_2242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(276), ack => WPIPE_Block2_start_1035_inst_req_0); -- 
    -- CP-element group 277:  transition  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1035_Update/req
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1035_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1035_Sample/ack
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1035_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1035_update_start_
      -- CP-element group 277: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1035_sample_completed_
      -- 
    ack_2243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1035_inst_ack_0, ack => convTranspose_CP_39_elements(277)); -- 
    req_2247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(277), ack => WPIPE_Block2_start_1035_inst_req_1); -- 
    -- CP-element group 278:  transition  input  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (6) 
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1038_Sample/req
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1038_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1038_sample_start_
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1035_Update/ack
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1035_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1035_update_completed_
      -- 
    ack_2248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1035_inst_ack_1, ack => convTranspose_CP_39_elements(278)); -- 
    req_2256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(278), ack => WPIPE_Block2_start_1038_inst_req_0); -- 
    -- CP-element group 279:  transition  input  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (6) 
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1038_Sample/ack
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1038_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1038_Update/req
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1038_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1038_update_start_
      -- CP-element group 279: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1038_sample_completed_
      -- 
    ack_2257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1038_inst_ack_0, ack => convTranspose_CP_39_elements(279)); -- 
    req_2261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(279), ack => WPIPE_Block2_start_1038_inst_req_1); -- 
    -- CP-element group 280:  transition  input  output  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (6) 
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1038_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1041_sample_start_
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1041_Sample/$entry
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1038_Update/ack
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1041_Sample/req
      -- CP-element group 280: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1038_update_completed_
      -- 
    ack_2262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1038_inst_ack_1, ack => convTranspose_CP_39_elements(280)); -- 
    req_2270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(280), ack => WPIPE_Block2_start_1041_inst_req_0); -- 
    -- CP-element group 281:  transition  input  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281:  members (6) 
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1041_update_start_
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1041_sample_completed_
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1041_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1041_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1041_Sample/ack
      -- CP-element group 281: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1041_Update/req
      -- 
    ack_2271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1041_inst_ack_0, ack => convTranspose_CP_39_elements(281)); -- 
    req_2275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(281), ack => WPIPE_Block2_start_1041_inst_req_1); -- 
    -- CP-element group 282:  transition  input  output  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (6) 
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1041_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1044_Sample/req
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1044_Sample/$entry
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1044_sample_start_
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1041_Update/ack
      -- CP-element group 282: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1041_Update/$exit
      -- 
    ack_2276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1041_inst_ack_1, ack => convTranspose_CP_39_elements(282)); -- 
    req_2284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(282), ack => WPIPE_Block2_start_1044_inst_req_0); -- 
    -- CP-element group 283:  transition  input  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (6) 
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1044_Update/req
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1044_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1044_Sample/ack
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1044_Sample/$exit
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1044_update_start_
      -- CP-element group 283: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1044_sample_completed_
      -- 
    ack_2285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1044_inst_ack_0, ack => convTranspose_CP_39_elements(283)); -- 
    req_2289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(283), ack => WPIPE_Block2_start_1044_inst_req_1); -- 
    -- CP-element group 284:  transition  input  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	319 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1044_Update/ack
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1044_Update/$exit
      -- CP-element group 284: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1044_update_completed_
      -- 
    ack_2290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1044_inst_ack_1, ack => convTranspose_CP_39_elements(284)); -- 
    -- CP-element group 285:  transition  input  output  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	398 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	286 
    -- CP-element group 285:  members (6) 
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1047_Update/req
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1047_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1047_Sample/ack
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1047_Sample/$exit
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1047_update_start_
      -- CP-element group 285: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1047_sample_completed_
      -- 
    ack_2299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1047_inst_ack_0, ack => convTranspose_CP_39_elements(285)); -- 
    req_2303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(285), ack => WPIPE_Block3_start_1047_inst_req_1); -- 
    -- CP-element group 286:  transition  input  output  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	285 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (6) 
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1050_Sample/$entry
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1050_sample_start_
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1050_Sample/req
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1047_Update/ack
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1047_Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1047_update_completed_
      -- 
    ack_2304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1047_inst_ack_1, ack => convTranspose_CP_39_elements(286)); -- 
    req_2312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(286), ack => WPIPE_Block3_start_1050_inst_req_0); -- 
    -- CP-element group 287:  transition  input  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (6) 
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1050_Sample/$exit
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1050_sample_completed_
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1050_Sample/ack
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1050_update_start_
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1050_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1050_Update/req
      -- 
    ack_2313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1050_inst_ack_0, ack => convTranspose_CP_39_elements(287)); -- 
    req_2317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(287), ack => WPIPE_Block3_start_1050_inst_req_1); -- 
    -- CP-element group 288:  transition  input  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (6) 
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1050_Update/$exit
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1050_Update/ack
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1050_update_completed_
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1053_Sample/req
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1053_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1053_sample_start_
      -- 
    ack_2318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1050_inst_ack_1, ack => convTranspose_CP_39_elements(288)); -- 
    req_2326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(288), ack => WPIPE_Block3_start_1053_inst_req_0); -- 
    -- CP-element group 289:  transition  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (6) 
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1053_Update/req
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1053_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1053_Sample/ack
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1053_Sample/$exit
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1053_update_start_
      -- CP-element group 289: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1053_sample_completed_
      -- 
    ack_2327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1053_inst_ack_0, ack => convTranspose_CP_39_elements(289)); -- 
    req_2331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(289), ack => WPIPE_Block3_start_1053_inst_req_1); -- 
    -- CP-element group 290:  transition  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (6) 
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1056_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1056_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1053_Update/ack
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1053_Update/$exit
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1053_update_completed_
      -- CP-element group 290: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1056_Sample/req
      -- 
    ack_2332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1053_inst_ack_1, ack => convTranspose_CP_39_elements(290)); -- 
    req_2340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(290), ack => WPIPE_Block3_start_1056_inst_req_0); -- 
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1056_sample_completed_
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1056_update_start_
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1056_Update/req
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1056_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1056_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1056_Sample/$exit
      -- 
    ack_2341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1056_inst_ack_0, ack => convTranspose_CP_39_elements(291)); -- 
    req_2345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(291), ack => WPIPE_Block3_start_1056_inst_req_1); -- 
    -- CP-element group 292:  transition  input  output  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (6) 
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1059_sample_start_
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1059_Sample/req
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1056_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1059_Sample/$entry
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1056_Update/ack
      -- CP-element group 292: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1056_Update/$exit
      -- 
    ack_2346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1056_inst_ack_1, ack => convTranspose_CP_39_elements(292)); -- 
    req_2354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(292), ack => WPIPE_Block3_start_1059_inst_req_0); -- 
    -- CP-element group 293:  transition  input  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1059_sample_completed_
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1059_update_start_
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1059_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1059_Sample/ack
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1059_Update/req
      -- CP-element group 293: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1059_Update/$entry
      -- 
    ack_2355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1059_inst_ack_0, ack => convTranspose_CP_39_elements(293)); -- 
    req_2359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(293), ack => WPIPE_Block3_start_1059_inst_req_1); -- 
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1059_update_completed_
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1059_Update/ack
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1062_Sample/req
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1062_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1059_Update/$exit
      -- CP-element group 294: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1062_sample_start_
      -- 
    ack_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1059_inst_ack_1, ack => convTranspose_CP_39_elements(294)); -- 
    req_2368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(294), ack => WPIPE_Block3_start_1062_inst_req_0); -- 
    -- CP-element group 295:  transition  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (6) 
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1062_Update/req
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1062_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1062_Sample/ack
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1062_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1062_update_start_
      -- CP-element group 295: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1062_sample_completed_
      -- 
    ack_2369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1062_inst_ack_0, ack => convTranspose_CP_39_elements(295)); -- 
    req_2373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(295), ack => WPIPE_Block3_start_1062_inst_req_1); -- 
    -- CP-element group 296:  transition  input  output  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296:  members (6) 
      -- CP-element group 296: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1062_Update/ack
      -- CP-element group 296: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1065_sample_start_
      -- CP-element group 296: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1062_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1062_update_completed_
      -- CP-element group 296: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1065_Sample/req
      -- CP-element group 296: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1065_Sample/$entry
      -- 
    ack_2374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1062_inst_ack_1, ack => convTranspose_CP_39_elements(296)); -- 
    req_2382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(296), ack => WPIPE_Block3_start_1065_inst_req_0); -- 
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1065_Update/req
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1065_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1065_Sample/ack
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1065_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1065_update_start_
      -- CP-element group 297: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1065_sample_completed_
      -- 
    ack_2383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1065_inst_ack_0, ack => convTranspose_CP_39_elements(297)); -- 
    req_2387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(297), ack => WPIPE_Block3_start_1065_inst_req_1); -- 
    -- CP-element group 298:  transition  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (6) 
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1068_sample_start_
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1065_Update/ack
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1068_Sample/req
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1068_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1065_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1065_update_completed_
      -- 
    ack_2388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1065_inst_ack_1, ack => convTranspose_CP_39_elements(298)); -- 
    req_2396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(298), ack => WPIPE_Block3_start_1068_inst_req_0); -- 
    -- CP-element group 299:  transition  input  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1068_Update/req
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1068_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1068_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1068_Sample/ack
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1068_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1068_update_start_
      -- 
    ack_2397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1068_inst_ack_0, ack => convTranspose_CP_39_elements(299)); -- 
    req_2401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(299), ack => WPIPE_Block3_start_1068_inst_req_1); -- 
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1068_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1071_Sample/req
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1071_Sample/$entry
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1068_Update/ack
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1068_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1071_sample_start_
      -- 
    ack_2402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1068_inst_ack_1, ack => convTranspose_CP_39_elements(300)); -- 
    req_2410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(300), ack => WPIPE_Block3_start_1071_inst_req_0); -- 
    -- CP-element group 301:  transition  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (6) 
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1071_Sample/ack
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1071_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1071_Update/req
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1071_Sample/$exit
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1071_update_start_
      -- CP-element group 301: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1071_sample_completed_
      -- 
    ack_2411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1071_inst_ack_0, ack => convTranspose_CP_39_elements(301)); -- 
    req_2415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(301), ack => WPIPE_Block3_start_1071_inst_req_1); -- 
    -- CP-element group 302:  transition  input  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (6) 
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1071_Update/$exit
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1074_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1071_Update/ack
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1071_update_completed_
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1074_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1074_Sample/req
      -- 
    ack_2416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1071_inst_ack_1, ack => convTranspose_CP_39_elements(302)); -- 
    req_2424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(302), ack => WPIPE_Block3_start_1074_inst_req_0); -- 
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1074_update_start_
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1074_Update/req
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1074_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1074_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1074_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1074_Sample/$exit
      -- 
    ack_2425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1074_inst_ack_0, ack => convTranspose_CP_39_elements(303)); -- 
    req_2429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(303), ack => WPIPE_Block3_start_1074_inst_req_1); -- 
    -- CP-element group 304:  transition  input  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (6) 
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1074_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1077_Sample/$entry
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1074_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1074_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1077_Sample/req
      -- CP-element group 304: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1077_sample_start_
      -- 
    ack_2430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1074_inst_ack_1, ack => convTranspose_CP_39_elements(304)); -- 
    req_2438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(304), ack => WPIPE_Block3_start_1077_inst_req_0); -- 
    -- CP-element group 305:  transition  input  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305:  members (6) 
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1077_Update/$entry
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1077_update_start_
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1077_sample_completed_
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1077_Update/req
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1077_Sample/$exit
      -- CP-element group 305: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1077_Sample/ack
      -- 
    ack_2439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1077_inst_ack_0, ack => convTranspose_CP_39_elements(305)); -- 
    req_2443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(305), ack => WPIPE_Block3_start_1077_inst_req_1); -- 
    -- CP-element group 306:  transition  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (6) 
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1077_update_completed_
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1077_Update/ack
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1077_Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1080_sample_start_
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1080_Sample/$entry
      -- CP-element group 306: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1080_Sample/req
      -- 
    ack_2444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1077_inst_ack_1, ack => convTranspose_CP_39_elements(306)); -- 
    req_2452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(306), ack => WPIPE_Block3_start_1080_inst_req_0); -- 
    -- CP-element group 307:  transition  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1080_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1080_update_start_
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1080_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1080_Sample/ack
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1080_Update/$entry
      -- CP-element group 307: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1080_Update/req
      -- 
    ack_2453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1080_inst_ack_0, ack => convTranspose_CP_39_elements(307)); -- 
    req_2457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(307), ack => WPIPE_Block3_start_1080_inst_req_1); -- 
    -- CP-element group 308:  transition  input  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (6) 
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1080_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1080_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1080_Update/ack
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1083_sample_start_
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1083_Sample/$entry
      -- CP-element group 308: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1083_Sample/req
      -- 
    ack_2458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1080_inst_ack_1, ack => convTranspose_CP_39_elements(308)); -- 
    req_2466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(308), ack => WPIPE_Block3_start_1083_inst_req_0); -- 
    -- CP-element group 309:  transition  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (6) 
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1083_sample_completed_
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1083_update_start_
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1083_Sample/$exit
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1083_Sample/ack
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1083_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1083_Update/req
      -- 
    ack_2467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1083_inst_ack_0, ack => convTranspose_CP_39_elements(309)); -- 
    req_2471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(309), ack => WPIPE_Block3_start_1083_inst_req_1); -- 
    -- CP-element group 310:  transition  input  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	319 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1083_update_completed_
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1083_Update/$exit
      -- CP-element group 310: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1083_Update/ack
      -- 
    ack_2472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1083_inst_ack_1, ack => convTranspose_CP_39_elements(310)); -- 
    -- CP-element group 311:  transition  input  output  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	398 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (6) 
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block0_done_1087_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block0_done_1087_update_start_
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block0_done_1087_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block0_done_1087_Sample/ra
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block0_done_1087_Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block0_done_1087_Update/cr
      -- 
    ra_2481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1087_inst_ack_0, ack => convTranspose_CP_39_elements(311)); -- 
    cr_2485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(311), ack => RPIPE_Block0_done_1087_inst_req_1); -- 
    -- CP-element group 312:  transition  input  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	319 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block0_done_1087_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block0_done_1087_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block0_done_1087_Update/ca
      -- 
    ca_2486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1087_inst_ack_1, ack => convTranspose_CP_39_elements(312)); -- 
    -- CP-element group 313:  transition  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	398 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (6) 
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block1_done_1090_sample_completed_
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block1_done_1090_update_start_
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block1_done_1090_Sample/$exit
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block1_done_1090_Sample/ra
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block1_done_1090_Update/$entry
      -- CP-element group 313: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block1_done_1090_Update/cr
      -- 
    ra_2495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1090_inst_ack_0, ack => convTranspose_CP_39_elements(313)); -- 
    cr_2499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(313), ack => RPIPE_Block1_done_1090_inst_req_1); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	319 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block1_done_1090_update_completed_
      -- CP-element group 314: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block1_done_1090_Update/$exit
      -- CP-element group 314: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block1_done_1090_Update/ca
      -- 
    ca_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1090_inst_ack_1, ack => convTranspose_CP_39_elements(314)); -- 
    -- CP-element group 315:  transition  input  output  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	398 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	316 
    -- CP-element group 315:  members (6) 
      -- CP-element group 315: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block2_done_1093_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block2_done_1093_update_start_
      -- CP-element group 315: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block2_done_1093_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block2_done_1093_Sample/ra
      -- CP-element group 315: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block2_done_1093_Update/$entry
      -- CP-element group 315: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block2_done_1093_Update/cr
      -- 
    ra_2509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1093_inst_ack_0, ack => convTranspose_CP_39_elements(315)); -- 
    cr_2513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(315), ack => RPIPE_Block2_done_1093_inst_req_1); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	315 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	319 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block2_done_1093_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block2_done_1093_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block2_done_1093_Update/ca
      -- 
    ca_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1093_inst_ack_1, ack => convTranspose_CP_39_elements(316)); -- 
    -- CP-element group 317:  transition  input  output  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	398 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (6) 
      -- CP-element group 317: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block3_done_1096_sample_completed_
      -- CP-element group 317: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block3_done_1096_update_start_
      -- CP-element group 317: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block3_done_1096_Sample/$exit
      -- CP-element group 317: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block3_done_1096_Sample/ra
      -- CP-element group 317: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block3_done_1096_Update/$entry
      -- CP-element group 317: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block3_done_1096_Update/cr
      -- 
    ra_2523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1096_inst_ack_0, ack => convTranspose_CP_39_elements(317)); -- 
    cr_2527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(317), ack => RPIPE_Block3_done_1096_inst_req_1); -- 
    -- CP-element group 318:  transition  input  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (3) 
      -- CP-element group 318: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block3_done_1096_update_completed_
      -- CP-element group 318: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block3_done_1096_Update/$exit
      -- CP-element group 318: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block3_done_1096_Update/ca
      -- 
    ca_2528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1096_inst_ack_1, ack => convTranspose_CP_39_elements(318)); -- 
    -- CP-element group 319:  join  fork  transition  place  output  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	206 
    -- CP-element group 319: 	232 
    -- CP-element group 319: 	258 
    -- CP-element group 319: 	284 
    -- CP-element group 319: 	310 
    -- CP-element group 319: 	312 
    -- CP-element group 319: 	314 
    -- CP-element group 319: 	316 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	320 
    -- CP-element group 319: 	321 
    -- CP-element group 319: 	323 
    -- CP-element group 319:  members (13) 
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097__exit__
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113__entry__
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/$exit
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/$entry
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/call_stmt_1100_sample_start_
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/call_stmt_1100_update_start_
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/call_stmt_1100_Sample/$entry
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/call_stmt_1100_Sample/crr
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/call_stmt_1100_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/call_stmt_1100_Update/ccr
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/type_cast_1104_update_start_
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/type_cast_1104_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/type_cast_1104_Update/cr
      -- 
    crr_2539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(319), ack => call_stmt_1100_call_req_0); -- 
    ccr_2544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(319), ack => call_stmt_1100_call_req_1); -- 
    cr_2558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(319), ack => type_cast_1104_inst_req_1); -- 
    convTranspose_cp_element_group_319: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_319"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(206) & convTranspose_CP_39_elements(232) & convTranspose_CP_39_elements(258) & convTranspose_CP_39_elements(284) & convTranspose_CP_39_elements(310) & convTranspose_CP_39_elements(312) & convTranspose_CP_39_elements(314) & convTranspose_CP_39_elements(316) & convTranspose_CP_39_elements(318);
      gj_convTranspose_cp_element_group_319 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(319), clk => clk, reset => reset); --
    end block;
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	319 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/call_stmt_1100_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/call_stmt_1100_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/call_stmt_1100_Sample/cra
      -- 
    cra_2540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1100_call_ack_0, ack => convTranspose_CP_39_elements(320)); -- 
    -- CP-element group 321:  transition  input  output  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	319 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (6) 
      -- CP-element group 321: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/call_stmt_1100_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/call_stmt_1100_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/call_stmt_1100_Update/cca
      -- CP-element group 321: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/type_cast_1104_sample_start_
      -- CP-element group 321: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/type_cast_1104_Sample/$entry
      -- CP-element group 321: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/type_cast_1104_Sample/rr
      -- 
    cca_2545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1100_call_ack_1, ack => convTranspose_CP_39_elements(321)); -- 
    rr_2553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(321), ack => type_cast_1104_inst_req_0); -- 
    -- CP-element group 322:  transition  input  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/type_cast_1104_sample_completed_
      -- CP-element group 322: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/type_cast_1104_Sample/$exit
      -- CP-element group 322: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/type_cast_1104_Sample/ra
      -- 
    ra_2554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1104_inst_ack_0, ack => convTranspose_CP_39_elements(322)); -- 
    -- CP-element group 323:  transition  input  output  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	319 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (6) 
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/type_cast_1104_update_completed_
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/type_cast_1104_Update/$exit
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/type_cast_1104_Update/ca
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/WPIPE_elapsed_time_pipe_1111_sample_start_
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/WPIPE_elapsed_time_pipe_1111_Sample/$entry
      -- CP-element group 323: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/WPIPE_elapsed_time_pipe_1111_Sample/req
      -- 
    ca_2559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1104_inst_ack_1, ack => convTranspose_CP_39_elements(323)); -- 
    req_2567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(323), ack => WPIPE_elapsed_time_pipe_1111_inst_req_0); -- 
    -- CP-element group 324:  transition  input  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (6) 
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/WPIPE_elapsed_time_pipe_1111_sample_completed_
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/WPIPE_elapsed_time_pipe_1111_update_start_
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/WPIPE_elapsed_time_pipe_1111_Sample/$exit
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/WPIPE_elapsed_time_pipe_1111_Sample/ack
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/WPIPE_elapsed_time_pipe_1111_Update/$entry
      -- CP-element group 324: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/WPIPE_elapsed_time_pipe_1111_Update/req
      -- 
    ack_2568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1111_inst_ack_0, ack => convTranspose_CP_39_elements(324)); -- 
    req_2572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(324), ack => WPIPE_elapsed_time_pipe_1111_inst_req_1); -- 
    -- CP-element group 325:  branch  transition  place  input  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325: 	327 
    -- CP-element group 325:  members (13) 
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113__exit__
      -- CP-element group 325: 	 branch_block_stmt_32/if_stmt_1115__entry__
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/$exit
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/WPIPE_elapsed_time_pipe_1111_update_completed_
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/WPIPE_elapsed_time_pipe_1111_Update/$exit
      -- CP-element group 325: 	 branch_block_stmt_32/call_stmt_1100_to_assign_stmt_1113/WPIPE_elapsed_time_pipe_1111_Update/ack
      -- CP-element group 325: 	 branch_block_stmt_32/if_stmt_1115_dead_link/$entry
      -- CP-element group 325: 	 branch_block_stmt_32/if_stmt_1115_eval_test/$entry
      -- CP-element group 325: 	 branch_block_stmt_32/if_stmt_1115_eval_test/$exit
      -- CP-element group 325: 	 branch_block_stmt_32/if_stmt_1115_eval_test/branch_req
      -- CP-element group 325: 	 branch_block_stmt_32/R_cmp264479_1116_place
      -- CP-element group 325: 	 branch_block_stmt_32/if_stmt_1115_if_link/$entry
      -- CP-element group 325: 	 branch_block_stmt_32/if_stmt_1115_else_link/$entry
      -- 
    ack_2573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1111_inst_ack_1, ack => convTranspose_CP_39_elements(325)); -- 
    branch_req_2581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(325), ack => if_stmt_1115_branch_req_0); -- 
    -- CP-element group 326:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	328 
    -- CP-element group 326: 	329 
    -- CP-element group 326:  members (18) 
      -- CP-element group 326: 	 branch_block_stmt_32/merge_stmt_1121__exit__
      -- CP-element group 326: 	 branch_block_stmt_32/assign_stmt_1127_to_assign_stmt_1156__entry__
      -- CP-element group 326: 	 branch_block_stmt_32/merge_stmt_1121_PhiReqMerge
      -- CP-element group 326: 	 branch_block_stmt_32/merge_stmt_1121_PhiAck/dummy
      -- CP-element group 326: 	 branch_block_stmt_32/merge_stmt_1121_PhiAck/$exit
      -- CP-element group 326: 	 branch_block_stmt_32/merge_stmt_1121_PhiAck/$entry
      -- CP-element group 326: 	 branch_block_stmt_32/forx_xend273_bbx_xnph_PhiReq/$exit
      -- CP-element group 326: 	 branch_block_stmt_32/forx_xend273_bbx_xnph_PhiReq/$entry
      -- CP-element group 326: 	 branch_block_stmt_32/if_stmt_1115_if_link/$exit
      -- CP-element group 326: 	 branch_block_stmt_32/if_stmt_1115_if_link/if_choice_transition
      -- CP-element group 326: 	 branch_block_stmt_32/forx_xend273_bbx_xnph
      -- CP-element group 326: 	 branch_block_stmt_32/assign_stmt_1127_to_assign_stmt_1156/$entry
      -- CP-element group 326: 	 branch_block_stmt_32/assign_stmt_1127_to_assign_stmt_1156/type_cast_1142_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_32/assign_stmt_1127_to_assign_stmt_1156/type_cast_1142_update_start_
      -- CP-element group 326: 	 branch_block_stmt_32/assign_stmt_1127_to_assign_stmt_1156/type_cast_1142_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_32/assign_stmt_1127_to_assign_stmt_1156/type_cast_1142_Sample/rr
      -- CP-element group 326: 	 branch_block_stmt_32/assign_stmt_1127_to_assign_stmt_1156/type_cast_1142_Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_32/assign_stmt_1127_to_assign_stmt_1156/type_cast_1142_Update/cr
      -- 
    if_choice_transition_2586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1115_branch_ack_1, ack => convTranspose_CP_39_elements(326)); -- 
    rr_2603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(326), ack => type_cast_1142_inst_req_0); -- 
    cr_2608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(326), ack => type_cast_1142_inst_req_1); -- 
    -- CP-element group 327:  transition  place  input  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	325 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	405 
    -- CP-element group 327:  members (5) 
      -- CP-element group 327: 	 branch_block_stmt_32/if_stmt_1115_else_link/$exit
      -- CP-element group 327: 	 branch_block_stmt_32/if_stmt_1115_else_link/else_choice_transition
      -- CP-element group 327: 	 branch_block_stmt_32/forx_xend273_forx_xend474
      -- CP-element group 327: 	 branch_block_stmt_32/forx_xend273_forx_xend474_PhiReq/$exit
      -- CP-element group 327: 	 branch_block_stmt_32/forx_xend273_forx_xend474_PhiReq/$entry
      -- 
    else_choice_transition_2590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1115_branch_ack_0, ack => convTranspose_CP_39_elements(327)); -- 
    -- CP-element group 328:  transition  input  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	326 
    -- CP-element group 328: successors 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 branch_block_stmt_32/assign_stmt_1127_to_assign_stmt_1156/type_cast_1142_sample_completed_
      -- CP-element group 328: 	 branch_block_stmt_32/assign_stmt_1127_to_assign_stmt_1156/type_cast_1142_Sample/$exit
      -- CP-element group 328: 	 branch_block_stmt_32/assign_stmt_1127_to_assign_stmt_1156/type_cast_1142_Sample/ra
      -- 
    ra_2604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1142_inst_ack_0, ack => convTranspose_CP_39_elements(328)); -- 
    -- CP-element group 329:  transition  place  input  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	326 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	399 
    -- CP-element group 329:  members (9) 
      -- CP-element group 329: 	 branch_block_stmt_32/assign_stmt_1127_to_assign_stmt_1156__exit__
      -- CP-element group 329: 	 branch_block_stmt_32/bbx_xnph_forx_xbody402
      -- CP-element group 329: 	 branch_block_stmt_32/bbx_xnph_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_sources/$entry
      -- CP-element group 329: 	 branch_block_stmt_32/bbx_xnph_forx_xbody402_PhiReq/phi_stmt_1159/$entry
      -- CP-element group 329: 	 branch_block_stmt_32/bbx_xnph_forx_xbody402_PhiReq/$entry
      -- CP-element group 329: 	 branch_block_stmt_32/assign_stmt_1127_to_assign_stmt_1156/$exit
      -- CP-element group 329: 	 branch_block_stmt_32/assign_stmt_1127_to_assign_stmt_1156/type_cast_1142_update_completed_
      -- CP-element group 329: 	 branch_block_stmt_32/assign_stmt_1127_to_assign_stmt_1156/type_cast_1142_Update/$exit
      -- CP-element group 329: 	 branch_block_stmt_32/assign_stmt_1127_to_assign_stmt_1156/type_cast_1142_Update/ca
      -- 
    ca_2609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1142_inst_ack_1, ack => convTranspose_CP_39_elements(329)); -- 
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	404 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	375 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_final_index_sum_regn_sample_complete
      -- CP-element group 330: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_final_index_sum_regn_Sample/$exit
      -- CP-element group 330: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_final_index_sum_regn_Sample/ack
      -- 
    ack_2638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1171_index_offset_ack_0, ack => convTranspose_CP_39_elements(330)); -- 
    -- CP-element group 331:  transition  input  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	404 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331:  members (11) 
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/addr_of_1172_sample_start_
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_root_address_calculated
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_offset_calculated
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_final_index_sum_regn_Update/$exit
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_final_index_sum_regn_Update/ack
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_base_plus_offset/$entry
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_base_plus_offset/$exit
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_base_plus_offset/sum_rename_req
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_base_plus_offset/sum_rename_ack
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/addr_of_1172_request/$entry
      -- CP-element group 331: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/addr_of_1172_request/req
      -- 
    ack_2643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1171_index_offset_ack_1, ack => convTranspose_CP_39_elements(331)); -- 
    req_2652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(331), ack => addr_of_1172_final_reg_req_0); -- 
    -- CP-element group 332:  transition  input  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/addr_of_1172_sample_completed_
      -- CP-element group 332: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/addr_of_1172_request/$exit
      -- CP-element group 332: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/addr_of_1172_request/ack
      -- 
    ack_2653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1172_final_reg_ack_0, ack => convTranspose_CP_39_elements(332)); -- 
    -- CP-element group 333:  join  fork  transition  input  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	404 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (24) 
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/addr_of_1172_update_completed_
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/addr_of_1172_complete/$exit
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/addr_of_1172_complete/ack
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_sample_start_
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_base_address_calculated
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_word_address_calculated
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_root_address_calculated
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_base_address_resized
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_base_addr_resize/$entry
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_base_addr_resize/$exit
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_base_addr_resize/base_resize_req
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_base_addr_resize/base_resize_ack
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_base_plus_offset/$entry
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_base_plus_offset/$exit
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_base_plus_offset/sum_rename_req
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_base_plus_offset/sum_rename_ack
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_word_addrgen/$entry
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_word_addrgen/$exit
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_word_addrgen/root_register_req
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_word_addrgen/root_register_ack
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Sample/$entry
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Sample/word_access_start/$entry
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Sample/word_access_start/word_0/$entry
      -- CP-element group 333: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Sample/word_access_start/word_0/rr
      -- 
    ack_2658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1172_final_reg_ack_1, ack => convTranspose_CP_39_elements(333)); -- 
    rr_2691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(333), ack => ptr_deref_1176_load_0_req_0); -- 
    -- CP-element group 334:  transition  input  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334:  members (5) 
      -- CP-element group 334: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_sample_completed_
      -- CP-element group 334: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Sample/$exit
      -- CP-element group 334: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Sample/word_access_start/$exit
      -- CP-element group 334: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Sample/word_access_start/word_0/$exit
      -- CP-element group 334: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Sample/word_access_start/word_0/ra
      -- 
    ra_2692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1176_load_0_ack_0, ack => convTranspose_CP_39_elements(334)); -- 
    -- CP-element group 335:  fork  transition  input  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	404 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	336 
    -- CP-element group 335: 	338 
    -- CP-element group 335: 	340 
    -- CP-element group 335: 	342 
    -- CP-element group 335: 	344 
    -- CP-element group 335: 	346 
    -- CP-element group 335: 	348 
    -- CP-element group 335: 	350 
    -- CP-element group 335:  members (33) 
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_update_completed_
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Update/$exit
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Update/word_access_complete/$exit
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Update/word_access_complete/word_0/$exit
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Update/word_access_complete/word_0/ca
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Update/ptr_deref_1176_Merge/$entry
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Update/ptr_deref_1176_Merge/$exit
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Update/ptr_deref_1176_Merge/merge_req
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Update/ptr_deref_1176_Merge/merge_ack
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1180_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1180_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1180_Sample/rr
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1190_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1190_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1190_Sample/rr
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1200_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1200_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1200_Sample/rr
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1210_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1210_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1210_Sample/rr
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1220_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1220_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1220_Sample/rr
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1230_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1230_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1230_Sample/rr
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1240_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1240_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1240_Sample/rr
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1250_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1250_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1250_Sample/rr
      -- 
    ca_2703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1176_load_0_ack_1, ack => convTranspose_CP_39_elements(335)); -- 
    rr_2716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(335), ack => type_cast_1180_inst_req_0); -- 
    rr_2730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(335), ack => type_cast_1190_inst_req_0); -- 
    rr_2744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(335), ack => type_cast_1200_inst_req_0); -- 
    rr_2758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(335), ack => type_cast_1210_inst_req_0); -- 
    rr_2772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(335), ack => type_cast_1220_inst_req_0); -- 
    rr_2786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(335), ack => type_cast_1230_inst_req_0); -- 
    rr_2800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(335), ack => type_cast_1240_inst_req_0); -- 
    rr_2814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(335), ack => type_cast_1250_inst_req_0); -- 
    -- CP-element group 336:  transition  input  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	335 
    -- CP-element group 336: successors 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1180_sample_completed_
      -- CP-element group 336: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1180_Sample/$exit
      -- CP-element group 336: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1180_Sample/ra
      -- 
    ra_2717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1180_inst_ack_0, ack => convTranspose_CP_39_elements(336)); -- 
    -- CP-element group 337:  transition  input  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	404 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	372 
    -- CP-element group 337:  members (3) 
      -- CP-element group 337: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1180_update_completed_
      -- CP-element group 337: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1180_Update/$exit
      -- CP-element group 337: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1180_Update/ca
      -- 
    ca_2722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1180_inst_ack_1, ack => convTranspose_CP_39_elements(337)); -- 
    -- CP-element group 338:  transition  input  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	335 
    -- CP-element group 338: successors 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1190_sample_completed_
      -- CP-element group 338: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1190_Sample/$exit
      -- CP-element group 338: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1190_Sample/ra
      -- 
    ra_2731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1190_inst_ack_0, ack => convTranspose_CP_39_elements(338)); -- 
    -- CP-element group 339:  transition  input  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	404 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	369 
    -- CP-element group 339:  members (3) 
      -- CP-element group 339: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1190_update_completed_
      -- CP-element group 339: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1190_Update/$exit
      -- CP-element group 339: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1190_Update/ca
      -- 
    ca_2736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1190_inst_ack_1, ack => convTranspose_CP_39_elements(339)); -- 
    -- CP-element group 340:  transition  input  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	335 
    -- CP-element group 340: successors 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1200_sample_completed_
      -- CP-element group 340: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1200_Sample/$exit
      -- CP-element group 340: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1200_Sample/ra
      -- 
    ra_2745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1200_inst_ack_0, ack => convTranspose_CP_39_elements(340)); -- 
    -- CP-element group 341:  transition  input  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	404 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	366 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1200_update_completed_
      -- CP-element group 341: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1200_Update/$exit
      -- CP-element group 341: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1200_Update/ca
      -- 
    ca_2750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1200_inst_ack_1, ack => convTranspose_CP_39_elements(341)); -- 
    -- CP-element group 342:  transition  input  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	335 
    -- CP-element group 342: successors 
    -- CP-element group 342:  members (3) 
      -- CP-element group 342: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1210_sample_completed_
      -- CP-element group 342: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1210_Sample/$exit
      -- CP-element group 342: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1210_Sample/ra
      -- 
    ra_2759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1210_inst_ack_0, ack => convTranspose_CP_39_elements(342)); -- 
    -- CP-element group 343:  transition  input  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	404 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	363 
    -- CP-element group 343:  members (3) 
      -- CP-element group 343: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1210_update_completed_
      -- CP-element group 343: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1210_Update/$exit
      -- CP-element group 343: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1210_Update/ca
      -- 
    ca_2764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1210_inst_ack_1, ack => convTranspose_CP_39_elements(343)); -- 
    -- CP-element group 344:  transition  input  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	335 
    -- CP-element group 344: successors 
    -- CP-element group 344:  members (3) 
      -- CP-element group 344: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1220_sample_completed_
      -- CP-element group 344: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1220_Sample/$exit
      -- CP-element group 344: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1220_Sample/ra
      -- 
    ra_2773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1220_inst_ack_0, ack => convTranspose_CP_39_elements(344)); -- 
    -- CP-element group 345:  transition  input  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	404 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	360 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1220_update_completed_
      -- CP-element group 345: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1220_Update/$exit
      -- CP-element group 345: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1220_Update/ca
      -- 
    ca_2778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1220_inst_ack_1, ack => convTranspose_CP_39_elements(345)); -- 
    -- CP-element group 346:  transition  input  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	335 
    -- CP-element group 346: successors 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1230_sample_completed_
      -- CP-element group 346: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1230_Sample/$exit
      -- CP-element group 346: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1230_Sample/ra
      -- 
    ra_2787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1230_inst_ack_0, ack => convTranspose_CP_39_elements(346)); -- 
    -- CP-element group 347:  transition  input  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	404 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	357 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1230_update_completed_
      -- CP-element group 347: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1230_Update/$exit
      -- CP-element group 347: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1230_Update/ca
      -- 
    ca_2792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1230_inst_ack_1, ack => convTranspose_CP_39_elements(347)); -- 
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	335 
    -- CP-element group 348: successors 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1240_sample_completed_
      -- CP-element group 348: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1240_Sample/$exit
      -- CP-element group 348: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1240_Sample/ra
      -- 
    ra_2801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1240_inst_ack_0, ack => convTranspose_CP_39_elements(348)); -- 
    -- CP-element group 349:  transition  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	404 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	354 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1240_update_completed_
      -- CP-element group 349: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1240_Update/$exit
      -- CP-element group 349: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1240_Update/ca
      -- 
    ca_2806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1240_inst_ack_1, ack => convTranspose_CP_39_elements(349)); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	335 
    -- CP-element group 350: successors 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1250_sample_completed_
      -- CP-element group 350: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1250_Sample/$exit
      -- CP-element group 350: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1250_Sample/ra
      -- 
    ra_2815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1250_inst_ack_0, ack => convTranspose_CP_39_elements(350)); -- 
    -- CP-element group 351:  transition  input  output  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	404 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (6) 
      -- CP-element group 351: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1250_update_completed_
      -- CP-element group 351: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1250_Update/$exit
      -- CP-element group 351: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1250_Update/ca
      -- CP-element group 351: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1252_sample_start_
      -- CP-element group 351: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1252_Sample/$entry
      -- CP-element group 351: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1252_Sample/req
      -- 
    ca_2820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1250_inst_ack_1, ack => convTranspose_CP_39_elements(351)); -- 
    req_2828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(351), ack => WPIPE_ConvTranspose_output_pipe_1252_inst_req_0); -- 
    -- CP-element group 352:  transition  input  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (6) 
      -- CP-element group 352: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1252_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1252_update_start_
      -- CP-element group 352: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1252_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1252_Sample/ack
      -- CP-element group 352: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1252_Update/$entry
      -- CP-element group 352: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1252_Update/req
      -- 
    ack_2829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1252_inst_ack_0, ack => convTranspose_CP_39_elements(352)); -- 
    req_2833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(352), ack => WPIPE_ConvTranspose_output_pipe_1252_inst_req_1); -- 
    -- CP-element group 353:  transition  input  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	354 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1252_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1252_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1252_Update/ack
      -- 
    ack_2834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1252_inst_ack_1, ack => convTranspose_CP_39_elements(353)); -- 
    -- CP-element group 354:  join  transition  output  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	349 
    -- CP-element group 354: 	353 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	355 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1255_sample_start_
      -- CP-element group 354: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1255_Sample/$entry
      -- CP-element group 354: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1255_Sample/req
      -- 
    req_2842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(354), ack => WPIPE_ConvTranspose_output_pipe_1255_inst_req_0); -- 
    convTranspose_cp_element_group_354: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_354"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(349) & convTranspose_CP_39_elements(353);
      gj_convTranspose_cp_element_group_354 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 355:  transition  input  output  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	354 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (6) 
      -- CP-element group 355: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1255_sample_completed_
      -- CP-element group 355: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1255_update_start_
      -- CP-element group 355: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1255_Sample/$exit
      -- CP-element group 355: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1255_Sample/ack
      -- CP-element group 355: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1255_Update/$entry
      -- CP-element group 355: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1255_Update/req
      -- 
    ack_2843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1255_inst_ack_0, ack => convTranspose_CP_39_elements(355)); -- 
    req_2847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(355), ack => WPIPE_ConvTranspose_output_pipe_1255_inst_req_1); -- 
    -- CP-element group 356:  transition  input  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1255_update_completed_
      -- CP-element group 356: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1255_Update/$exit
      -- CP-element group 356: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1255_Update/ack
      -- 
    ack_2848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1255_inst_ack_1, ack => convTranspose_CP_39_elements(356)); -- 
    -- CP-element group 357:  join  transition  output  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	347 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1258_sample_start_
      -- CP-element group 357: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1258_Sample/$entry
      -- CP-element group 357: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1258_Sample/req
      -- 
    req_2856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(357), ack => WPIPE_ConvTranspose_output_pipe_1258_inst_req_0); -- 
    convTranspose_cp_element_group_357: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_357"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(347) & convTranspose_CP_39_elements(356);
      gj_convTranspose_cp_element_group_357 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(357), clk => clk, reset => reset); --
    end block;
    -- CP-element group 358:  transition  input  output  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (6) 
      -- CP-element group 358: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1258_sample_completed_
      -- CP-element group 358: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1258_update_start_
      -- CP-element group 358: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1258_Sample/$exit
      -- CP-element group 358: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1258_Sample/ack
      -- CP-element group 358: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1258_Update/$entry
      -- CP-element group 358: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1258_Update/req
      -- 
    ack_2857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1258_inst_ack_0, ack => convTranspose_CP_39_elements(358)); -- 
    req_2861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(358), ack => WPIPE_ConvTranspose_output_pipe_1258_inst_req_1); -- 
    -- CP-element group 359:  transition  input  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	360 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1258_update_completed_
      -- CP-element group 359: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1258_Update/$exit
      -- CP-element group 359: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1258_Update/ack
      -- 
    ack_2862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1258_inst_ack_1, ack => convTranspose_CP_39_elements(359)); -- 
    -- CP-element group 360:  join  transition  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	345 
    -- CP-element group 360: 	359 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1261_sample_start_
      -- CP-element group 360: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1261_Sample/$entry
      -- CP-element group 360: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1261_Sample/req
      -- 
    req_2870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(360), ack => WPIPE_ConvTranspose_output_pipe_1261_inst_req_0); -- 
    convTranspose_cp_element_group_360: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_360"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(345) & convTranspose_CP_39_elements(359);
      gj_convTranspose_cp_element_group_360 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(360), clk => clk, reset => reset); --
    end block;
    -- CP-element group 361:  transition  input  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (6) 
      -- CP-element group 361: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1261_sample_completed_
      -- CP-element group 361: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1261_update_start_
      -- CP-element group 361: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1261_Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1261_Sample/ack
      -- CP-element group 361: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1261_Update/$entry
      -- CP-element group 361: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1261_Update/req
      -- 
    ack_2871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1261_inst_ack_0, ack => convTranspose_CP_39_elements(361)); -- 
    req_2875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(361), ack => WPIPE_ConvTranspose_output_pipe_1261_inst_req_1); -- 
    -- CP-element group 362:  transition  input  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	363 
    -- CP-element group 362:  members (3) 
      -- CP-element group 362: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1261_update_completed_
      -- CP-element group 362: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1261_Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1261_Update/ack
      -- 
    ack_2876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1261_inst_ack_1, ack => convTranspose_CP_39_elements(362)); -- 
    -- CP-element group 363:  join  transition  output  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	343 
    -- CP-element group 363: 	362 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (3) 
      -- CP-element group 363: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1264_sample_start_
      -- CP-element group 363: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1264_Sample/$entry
      -- CP-element group 363: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1264_Sample/req
      -- 
    req_2884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(363), ack => WPIPE_ConvTranspose_output_pipe_1264_inst_req_0); -- 
    convTranspose_cp_element_group_363: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_363"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(343) & convTranspose_CP_39_elements(362);
      gj_convTranspose_cp_element_group_363 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(363), clk => clk, reset => reset); --
    end block;
    -- CP-element group 364:  transition  input  output  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (6) 
      -- CP-element group 364: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1264_sample_completed_
      -- CP-element group 364: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1264_update_start_
      -- CP-element group 364: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1264_Sample/$exit
      -- CP-element group 364: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1264_Sample/ack
      -- CP-element group 364: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1264_Update/$entry
      -- CP-element group 364: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1264_Update/req
      -- 
    ack_2885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1264_inst_ack_0, ack => convTranspose_CP_39_elements(364)); -- 
    req_2889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(364), ack => WPIPE_ConvTranspose_output_pipe_1264_inst_req_1); -- 
    -- CP-element group 365:  transition  input  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (3) 
      -- CP-element group 365: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1264_update_completed_
      -- CP-element group 365: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1264_Update/$exit
      -- CP-element group 365: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1264_Update/ack
      -- 
    ack_2890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1264_inst_ack_1, ack => convTranspose_CP_39_elements(365)); -- 
    -- CP-element group 366:  join  transition  output  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	341 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	367 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1267_sample_start_
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1267_Sample/$entry
      -- CP-element group 366: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1267_Sample/req
      -- 
    req_2898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(366), ack => WPIPE_ConvTranspose_output_pipe_1267_inst_req_0); -- 
    convTranspose_cp_element_group_366: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_366"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(341) & convTranspose_CP_39_elements(365);
      gj_convTranspose_cp_element_group_366 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(366), clk => clk, reset => reset); --
    end block;
    -- CP-element group 367:  transition  input  output  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	366 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (6) 
      -- CP-element group 367: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1267_sample_completed_
      -- CP-element group 367: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1267_update_start_
      -- CP-element group 367: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1267_Sample/$exit
      -- CP-element group 367: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1267_Sample/ack
      -- CP-element group 367: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1267_Update/$entry
      -- CP-element group 367: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1267_Update/req
      -- 
    ack_2899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1267_inst_ack_0, ack => convTranspose_CP_39_elements(367)); -- 
    req_2903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(367), ack => WPIPE_ConvTranspose_output_pipe_1267_inst_req_1); -- 
    -- CP-element group 368:  transition  input  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	369 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1267_update_completed_
      -- CP-element group 368: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1267_Update/$exit
      -- CP-element group 368: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1267_Update/ack
      -- 
    ack_2904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1267_inst_ack_1, ack => convTranspose_CP_39_elements(368)); -- 
    -- CP-element group 369:  join  transition  output  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	339 
    -- CP-element group 369: 	368 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (3) 
      -- CP-element group 369: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1270_sample_start_
      -- CP-element group 369: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1270_Sample/$entry
      -- CP-element group 369: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1270_Sample/req
      -- 
    req_2912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(369), ack => WPIPE_ConvTranspose_output_pipe_1270_inst_req_0); -- 
    convTranspose_cp_element_group_369: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_369"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(339) & convTranspose_CP_39_elements(368);
      gj_convTranspose_cp_element_group_369 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(369), clk => clk, reset => reset); --
    end block;
    -- CP-element group 370:  transition  input  output  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370:  members (6) 
      -- CP-element group 370: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1270_sample_completed_
      -- CP-element group 370: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1270_update_start_
      -- CP-element group 370: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1270_Sample/$exit
      -- CP-element group 370: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1270_Sample/ack
      -- CP-element group 370: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1270_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1270_Update/req
      -- 
    ack_2913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1270_inst_ack_0, ack => convTranspose_CP_39_elements(370)); -- 
    req_2917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(370), ack => WPIPE_ConvTranspose_output_pipe_1270_inst_req_1); -- 
    -- CP-element group 371:  transition  input  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1270_update_completed_
      -- CP-element group 371: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1270_Update/$exit
      -- CP-element group 371: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1270_Update/ack
      -- 
    ack_2918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1270_inst_ack_1, ack => convTranspose_CP_39_elements(371)); -- 
    -- CP-element group 372:  join  transition  output  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	337 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1273_sample_start_
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1273_Sample/$entry
      -- CP-element group 372: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1273_Sample/req
      -- 
    req_2926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(372), ack => WPIPE_ConvTranspose_output_pipe_1273_inst_req_0); -- 
    convTranspose_cp_element_group_372: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_372"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(337) & convTranspose_CP_39_elements(371);
      gj_convTranspose_cp_element_group_372 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(372), clk => clk, reset => reset); --
    end block;
    -- CP-element group 373:  transition  input  output  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (6) 
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1273_sample_completed_
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1273_update_start_
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1273_Sample/$exit
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1273_Sample/ack
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1273_Update/$entry
      -- CP-element group 373: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1273_Update/req
      -- 
    ack_2927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1273_inst_ack_0, ack => convTranspose_CP_39_elements(373)); -- 
    req_2931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(373), ack => WPIPE_ConvTranspose_output_pipe_1273_inst_req_1); -- 
    -- CP-element group 374:  transition  input  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	375 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1273_update_completed_
      -- CP-element group 374: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1273_Update/$exit
      -- CP-element group 374: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/WPIPE_ConvTranspose_output_pipe_1273_Update/ack
      -- 
    ack_2932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1273_inst_ack_1, ack => convTranspose_CP_39_elements(374)); -- 
    -- CP-element group 375:  branch  join  transition  place  output  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	330 
    -- CP-element group 375: 	374 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	376 
    -- CP-element group 375: 	377 
    -- CP-element group 375:  members (10) 
      -- CP-element group 375: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286__exit__
      -- CP-element group 375: 	 branch_block_stmt_32/if_stmt_1287__entry__
      -- CP-element group 375: 	 branch_block_stmt_32/if_stmt_1287_else_link/$entry
      -- CP-element group 375: 	 branch_block_stmt_32/if_stmt_1287_if_link/$entry
      -- CP-element group 375: 	 branch_block_stmt_32/if_stmt_1287_eval_test/branch_req
      -- CP-element group 375: 	 branch_block_stmt_32/R_exitcond1_1288_place
      -- CP-element group 375: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/$exit
      -- CP-element group 375: 	 branch_block_stmt_32/if_stmt_1287_eval_test/$exit
      -- CP-element group 375: 	 branch_block_stmt_32/if_stmt_1287_eval_test/$entry
      -- CP-element group 375: 	 branch_block_stmt_32/if_stmt_1287_dead_link/$entry
      -- 
    branch_req_2940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(375), ack => if_stmt_1287_branch_req_0); -- 
    convTranspose_cp_element_group_375: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_375"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(330) & convTranspose_CP_39_elements(374);
      gj_convTranspose_cp_element_group_375 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(375), clk => clk, reset => reset); --
    end block;
    -- CP-element group 376:  merge  transition  place  input  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	375 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	405 
    -- CP-element group 376:  members (13) 
      -- CP-element group 376: 	 branch_block_stmt_32/merge_stmt_1293__exit__
      -- CP-element group 376: 	 branch_block_stmt_32/forx_xend474x_xloopexit_forx_xend474
      -- CP-element group 376: 	 branch_block_stmt_32/if_stmt_1287_if_link/$exit
      -- CP-element group 376: 	 branch_block_stmt_32/merge_stmt_1293_PhiReqMerge
      -- CP-element group 376: 	 branch_block_stmt_32/if_stmt_1287_if_link/if_choice_transition
      -- CP-element group 376: 	 branch_block_stmt_32/forx_xbody402_forx_xend474x_xloopexit
      -- CP-element group 376: 	 branch_block_stmt_32/forx_xend474x_xloopexit_forx_xend474_PhiReq/$exit
      -- CP-element group 376: 	 branch_block_stmt_32/forx_xend474x_xloopexit_forx_xend474_PhiReq/$entry
      -- CP-element group 376: 	 branch_block_stmt_32/merge_stmt_1293_PhiAck/dummy
      -- CP-element group 376: 	 branch_block_stmt_32/merge_stmt_1293_PhiAck/$exit
      -- CP-element group 376: 	 branch_block_stmt_32/merge_stmt_1293_PhiAck/$entry
      -- CP-element group 376: 	 branch_block_stmt_32/forx_xbody402_forx_xend474x_xloopexit_PhiReq/$exit
      -- CP-element group 376: 	 branch_block_stmt_32/forx_xbody402_forx_xend474x_xloopexit_PhiReq/$entry
      -- 
    if_choice_transition_2945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1287_branch_ack_1, ack => convTranspose_CP_39_elements(376)); -- 
    -- CP-element group 377:  fork  transition  place  input  output  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	375 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	400 
    -- CP-element group 377: 	401 
    -- CP-element group 377:  members (12) 
      -- CP-element group 377: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_sources/type_cast_1162/SplitProtocol/Sample/rr
      -- CP-element group 377: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_sources/type_cast_1162/SplitProtocol/Update/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_sources/type_cast_1162/SplitProtocol/Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_sources/type_cast_1162/SplitProtocol/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_sources/type_cast_1162/SplitProtocol/Update/cr
      -- CP-element group 377: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_sources/type_cast_1162/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/if_stmt_1287_else_link/$exit
      -- CP-element group 377: 	 branch_block_stmt_32/if_stmt_1287_else_link/else_choice_transition
      -- CP-element group 377: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_sources/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/phi_stmt_1159/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/$entry
      -- CP-element group 377: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402
      -- 
    else_choice_transition_2949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1287_branch_ack_0, ack => convTranspose_CP_39_elements(377)); -- 
    rr_3224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1162_inst_req_0); -- 
    cr_3229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(377), ack => type_cast_1162_inst_req_1); -- 
    -- CP-element group 378:  merge  branch  transition  place  output  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	144 
    -- CP-element group 378: 	99 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	100 
    -- CP-element group 378: 	101 
    -- CP-element group 378:  members (17) 
      -- CP-element group 378: 	 branch_block_stmt_32/merge_stmt_396__exit__
      -- CP-element group 378: 	 branch_block_stmt_32/assign_stmt_402__entry__
      -- CP-element group 378: 	 branch_block_stmt_32/assign_stmt_402__exit__
      -- CP-element group 378: 	 branch_block_stmt_32/if_stmt_403__entry__
      -- CP-element group 378: 	 branch_block_stmt_32/merge_stmt_396_PhiAck/dummy
      -- CP-element group 378: 	 branch_block_stmt_32/assign_stmt_402/$entry
      -- CP-element group 378: 	 branch_block_stmt_32/assign_stmt_402/$exit
      -- CP-element group 378: 	 branch_block_stmt_32/if_stmt_403_dead_link/$entry
      -- CP-element group 378: 	 branch_block_stmt_32/if_stmt_403_eval_test/$entry
      -- CP-element group 378: 	 branch_block_stmt_32/if_stmt_403_eval_test/$exit
      -- CP-element group 378: 	 branch_block_stmt_32/if_stmt_403_eval_test/branch_req
      -- CP-element group 378: 	 branch_block_stmt_32/R_cmp194483_404_place
      -- CP-element group 378: 	 branch_block_stmt_32/if_stmt_403_if_link/$entry
      -- CP-element group 378: 	 branch_block_stmt_32/if_stmt_403_else_link/$entry
      -- CP-element group 378: 	 branch_block_stmt_32/merge_stmt_396_PhiAck/$exit
      -- CP-element group 378: 	 branch_block_stmt_32/merge_stmt_396_PhiReqMerge
      -- CP-element group 378: 	 branch_block_stmt_32/merge_stmt_396_PhiAck/$entry
      -- 
    branch_req_827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(378), ack => if_stmt_403_branch_req_0); -- 
    convTranspose_CP_39_elements(378) <= OrReduce(convTranspose_CP_39_elements(144) & convTranspose_CP_39_elements(99));
    -- CP-element group 379:  transition  output  delay-element  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	103 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	383 
    -- CP-element group 379:  members (5) 
      -- CP-element group 379: 	 branch_block_stmt_32/bbx_xnph489_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_req
      -- CP-element group 379: 	 branch_block_stmt_32/bbx_xnph489_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_445_konst_delay_trans
      -- CP-element group 379: 	 branch_block_stmt_32/bbx_xnph489_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/$exit
      -- CP-element group 379: 	 branch_block_stmt_32/bbx_xnph489_forx_xbody_PhiReq/phi_stmt_441/$exit
      -- CP-element group 379: 	 branch_block_stmt_32/bbx_xnph489_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_441_req_2997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_441_req_2997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(379), ack => phi_stmt_441_req_0); -- 
    -- Element group convTranspose_CP_39_elements(379) is a control-delay.
    cp_element_379_delay: control_delay_element  generic map(name => " 379_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(103), ack => convTranspose_CP_39_elements(379), clk => clk, reset =>reset);
    -- CP-element group 380:  transition  input  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	145 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	382 
    -- CP-element group 380:  members (2) 
      -- CP-element group 380: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/Sample/$exit
      -- CP-element group 380: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/Sample/ra
      -- 
    ra_3017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_447_inst_ack_0, ack => convTranspose_CP_39_elements(380)); -- 
    -- CP-element group 381:  transition  input  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	145 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	382 
    -- CP-element group 381:  members (2) 
      -- CP-element group 381: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/Update/$exit
      -- CP-element group 381: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/Update/ca
      -- 
    ca_3022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_447_inst_ack_1, ack => convTranspose_CP_39_elements(381)); -- 
    -- CP-element group 382:  join  transition  output  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	380 
    -- CP-element group 382: 	381 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	383 
    -- CP-element group 382:  members (6) 
      -- CP-element group 382: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/$exit
      -- CP-element group 382: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/$exit
      -- CP-element group 382: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/SplitProtocol/$exit
      -- CP-element group 382: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_sources/type_cast_447/$exit
      -- CP-element group 382: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 382: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_441/phi_stmt_441_req
      -- 
    phi_stmt_441_req_3023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_441_req_3023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(382), ack => phi_stmt_441_req_1); -- 
    convTranspose_cp_element_group_382: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_382"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(380) & convTranspose_CP_39_elements(381);
      gj_convTranspose_cp_element_group_382 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(382), clk => clk, reset => reset); --
    end block;
    -- CP-element group 383:  merge  transition  place  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	379 
    -- CP-element group 383: 	382 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383:  members (2) 
      -- CP-element group 383: 	 branch_block_stmt_32/merge_stmt_440_PhiReqMerge
      -- CP-element group 383: 	 branch_block_stmt_32/merge_stmt_440_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(383) <= OrReduce(convTranspose_CP_39_elements(379) & convTranspose_CP_39_elements(382));
    -- CP-element group 384:  fork  transition  place  input  output  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	115 
    -- CP-element group 384: 	119 
    -- CP-element group 384: 	123 
    -- CP-element group 384: 	127 
    -- CP-element group 384: 	131 
    -- CP-element group 384: 	135 
    -- CP-element group 384: 	139 
    -- CP-element group 384: 	142 
    -- CP-element group 384: 	104 
    -- CP-element group 384: 	105 
    -- CP-element group 384: 	107 
    -- CP-element group 384: 	108 
    -- CP-element group 384: 	111 
    -- CP-element group 384:  members (56) 
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_492_update_start_
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_474_Update/cr
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Update/word_access_complete/word_0/cr
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_564_update_start_
      -- CP-element group 384: 	 branch_block_stmt_32/merge_stmt_440__exit__
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603__entry__
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_528_Update/cr
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_update_start_
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Update/word_access_complete/word_0/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Update/word_access_complete/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_528_update_start_
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/ptr_deref_590_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_582_Update/cr
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_582_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_492_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_564_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_582_update_start_
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_510_Update/cr
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_510_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_510_update_start_
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_546_Update/cr
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_546_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_492_Update/cr
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_564_Update/cr
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_528_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_474_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_546_update_start_
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/addr_of_454_update_start_
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_index_resized_1
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_index_scaled_1
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_index_computed_1
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_index_resize_1/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_index_resize_1/$exit
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_index_resize_1/index_resize_req
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_index_resize_1/index_resize_ack
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_index_scale_1/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_index_scale_1/$exit
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_index_scale_1/scale_rename_req
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_index_scale_1/scale_rename_ack
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_final_index_sum_regn_update_start
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_final_index_sum_regn_Sample/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_final_index_sum_regn_Sample/req
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_final_index_sum_regn_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/array_obj_ref_453_final_index_sum_regn_Update/req
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/addr_of_454_complete/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/addr_of_454_complete/req
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_457_sample_start_
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_457_Sample/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/RPIPE_ConvTranspose_input_pipe_457_Sample/rr
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_461_update_start_
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_461_Update/$entry
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_461_Update/cr
      -- CP-element group 384: 	 branch_block_stmt_32/assign_stmt_455_to_assign_stmt_603/type_cast_474_update_start_
      -- CP-element group 384: 	 branch_block_stmt_32/merge_stmt_440_PhiAck/phi_stmt_441_ack
      -- CP-element group 384: 	 branch_block_stmt_32/merge_stmt_440_PhiAck/$exit
      -- 
    phi_stmt_441_ack_3028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_441_ack_0, ack => convTranspose_CP_39_elements(384)); -- 
    cr_959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(384), ack => type_cast_474_inst_req_1); -- 
    cr_1177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(384), ack => ptr_deref_590_store_0_req_1); -- 
    cr_1043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(384), ack => type_cast_528_inst_req_1); -- 
    cr_1127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(384), ack => type_cast_582_inst_req_1); -- 
    cr_1015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(384), ack => type_cast_510_inst_req_1); -- 
    cr_1071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(384), ack => type_cast_546_inst_req_1); -- 
    cr_987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(384), ack => type_cast_492_inst_req_1); -- 
    cr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(384), ack => type_cast_564_inst_req_1); -- 
    req_883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(384), ack => array_obj_ref_453_index_offset_req_0); -- 
    req_888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(384), ack => array_obj_ref_453_index_offset_req_1); -- 
    req_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(384), ack => addr_of_454_final_reg_req_1); -- 
    rr_912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(384), ack => RPIPE_ConvTranspose_input_pipe_457_inst_req_0); -- 
    cr_931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(384), ack => type_cast_461_inst_req_1); -- 
    -- CP-element group 385:  transition  output  delay-element  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	147 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	389 
    -- CP-element group 385:  members (5) 
      -- CP-element group 385: 	 branch_block_stmt_32/bbx_xnph485_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_req
      -- CP-element group 385: 	 branch_block_stmt_32/bbx_xnph485_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_sources/type_cast_654_konst_delay_trans
      -- CP-element group 385: 	 branch_block_stmt_32/bbx_xnph485_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_sources/$exit
      -- CP-element group 385: 	 branch_block_stmt_32/bbx_xnph485_forx_xbody196_PhiReq/phi_stmt_648/$exit
      -- CP-element group 385: 	 branch_block_stmt_32/bbx_xnph485_forx_xbody196_PhiReq/$exit
      -- 
    phi_stmt_648_req_3051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_648_req_3051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(385), ack => phi_stmt_648_req_1); -- 
    -- Element group convTranspose_CP_39_elements(385) is a control-delay.
    cp_element_385_delay: control_delay_element  generic map(name => " 385_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(147), ack => convTranspose_CP_39_elements(385), clk => clk, reset =>reset);
    -- CP-element group 386:  transition  input  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	189 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	388 
    -- CP-element group 386:  members (2) 
      -- CP-element group 386: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_sources/type_cast_651/SplitProtocol/Sample/ra
      -- CP-element group 386: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_sources/type_cast_651/SplitProtocol/Sample/$exit
      -- 
    ra_3071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_651_inst_ack_0, ack => convTranspose_CP_39_elements(386)); -- 
    -- CP-element group 387:  transition  input  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	189 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	388 
    -- CP-element group 387:  members (2) 
      -- CP-element group 387: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_sources/type_cast_651/SplitProtocol/Update/ca
      -- CP-element group 387: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_sources/type_cast_651/SplitProtocol/Update/$exit
      -- 
    ca_3076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_651_inst_ack_1, ack => convTranspose_CP_39_elements(387)); -- 
    -- CP-element group 388:  join  transition  output  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	386 
    -- CP-element group 388: 	387 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	389 
    -- CP-element group 388:  members (6) 
      -- CP-element group 388: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_req
      -- CP-element group 388: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_sources/type_cast_651/SplitProtocol/$exit
      -- CP-element group 388: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_sources/type_cast_651/$exit
      -- CP-element group 388: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_648/phi_stmt_648_sources/$exit
      -- CP-element group 388: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/phi_stmt_648/$exit
      -- CP-element group 388: 	 branch_block_stmt_32/forx_xbody196_forx_xbody196_PhiReq/$exit
      -- 
    phi_stmt_648_req_3077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_648_req_3077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(388), ack => phi_stmt_648_req_0); -- 
    convTranspose_cp_element_group_388: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_388"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(386) & convTranspose_CP_39_elements(387);
      gj_convTranspose_cp_element_group_388 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(388), clk => clk, reset => reset); --
    end block;
    -- CP-element group 389:  merge  transition  place  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	385 
    -- CP-element group 389: 	388 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	390 
    -- CP-element group 389:  members (2) 
      -- CP-element group 389: 	 branch_block_stmt_32/merge_stmt_647_PhiReqMerge
      -- CP-element group 389: 	 branch_block_stmt_32/merge_stmt_647_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(389) <= OrReduce(convTranspose_CP_39_elements(385) & convTranspose_CP_39_elements(388));
    -- CP-element group 390:  fork  transition  place  input  output  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	389 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	148 
    -- CP-element group 390: 	149 
    -- CP-element group 390: 	151 
    -- CP-element group 390: 	152 
    -- CP-element group 390: 	155 
    -- CP-element group 390: 	159 
    -- CP-element group 390: 	163 
    -- CP-element group 390: 	167 
    -- CP-element group 390: 	171 
    -- CP-element group 390: 	175 
    -- CP-element group 390: 	179 
    -- CP-element group 390: 	183 
    -- CP-element group 390: 	186 
    -- CP-element group 390:  members (56) 
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_717_update_start_
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_735_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_735_Update/cr
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_668_update_start_
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_717_Update/cr
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_index_scaled_1
      -- CP-element group 390: 	 branch_block_stmt_32/merge_stmt_647__exit__
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810__entry__
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_index_resized_1
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_664_sample_start_
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_735_update_start_
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_681_Update/cr
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_681_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/addr_of_661_update_start_
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_final_index_sum_regn_Update/req
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_final_index_sum_regn_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_681_update_start_
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_final_index_sum_regn_Sample/req
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_699_Update/cr
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_index_resize_1/$exit
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_index_resize_1/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_699_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_664_Sample/rr
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_final_index_sum_regn_Sample/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/RPIPE_ConvTranspose_input_pipe_664_Sample/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_final_index_sum_regn_update_start
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/addr_of_661_complete/req
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_index_scale_1/scale_rename_ack
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_717_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_index_scale_1/scale_rename_req
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/addr_of_661_complete/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_index_scale_1/$exit
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_index_scale_1/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_668_Update/cr
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_index_resize_1/index_resize_ack
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_699_update_start_
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_668_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_index_resize_1/index_resize_req
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/array_obj_ref_660_index_computed_1
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_753_update_start_
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_753_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_753_Update/cr
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_771_update_start_
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_771_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_771_Update/cr
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_789_update_start_
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_789_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/type_cast_789_Update/cr
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_update_start_
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Update/word_access_complete/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Update/word_access_complete/word_0/$entry
      -- CP-element group 390: 	 branch_block_stmt_32/assign_stmt_662_to_assign_stmt_810/ptr_deref_797_Update/word_access_complete/word_0/cr
      -- CP-element group 390: 	 branch_block_stmt_32/merge_stmt_647_PhiAck/phi_stmt_648_ack
      -- CP-element group 390: 	 branch_block_stmt_32/merge_stmt_647_PhiAck/$exit
      -- 
    phi_stmt_648_ack_3082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_648_ack_0, ack => convTranspose_CP_39_elements(390)); -- 
    cr_1402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(390), ack => type_cast_735_inst_req_1); -- 
    cr_1374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(390), ack => type_cast_717_inst_req_1); -- 
    cr_1318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(390), ack => type_cast_681_inst_req_1); -- 
    req_1247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(390), ack => array_obj_ref_660_index_offset_req_1); -- 
    req_1242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(390), ack => array_obj_ref_660_index_offset_req_0); -- 
    cr_1346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(390), ack => type_cast_699_inst_req_1); -- 
    rr_1271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(390), ack => RPIPE_ConvTranspose_input_pipe_664_inst_req_0); -- 
    req_1262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(390), ack => addr_of_661_final_reg_req_1); -- 
    cr_1290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(390), ack => type_cast_668_inst_req_1); -- 
    cr_1430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(390), ack => type_cast_753_inst_req_1); -- 
    cr_1458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(390), ack => type_cast_771_inst_req_1); -- 
    cr_1486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(390), ack => type_cast_789_inst_req_1); -- 
    cr_1536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(390), ack => ptr_deref_797_store_0_req_1); -- 
    -- CP-element group 391:  merge  branch  transition  place  output  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	188 
    -- CP-element group 391: 	101 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	190 
    -- CP-element group 391: 	191 
    -- CP-element group 391:  members (17) 
      -- CP-element group 391: 	 branch_block_stmt_32/merge_stmt_819__exit__
      -- CP-element group 391: 	 branch_block_stmt_32/assign_stmt_824_to_assign_stmt_835__entry__
      -- CP-element group 391: 	 branch_block_stmt_32/assign_stmt_824_to_assign_stmt_835__exit__
      -- CP-element group 391: 	 branch_block_stmt_32/if_stmt_836__entry__
      -- CP-element group 391: 	 branch_block_stmt_32/merge_stmt_819_PhiReqMerge
      -- CP-element group 391: 	 branch_block_stmt_32/assign_stmt_824_to_assign_stmt_835/$entry
      -- CP-element group 391: 	 branch_block_stmt_32/assign_stmt_824_to_assign_stmt_835/$exit
      -- CP-element group 391: 	 branch_block_stmt_32/if_stmt_836_dead_link/$entry
      -- CP-element group 391: 	 branch_block_stmt_32/if_stmt_836_eval_test/$entry
      -- CP-element group 391: 	 branch_block_stmt_32/if_stmt_836_eval_test/$exit
      -- CP-element group 391: 	 branch_block_stmt_32/if_stmt_836_eval_test/branch_req
      -- CP-element group 391: 	 branch_block_stmt_32/R_cmp264479_837_place
      -- CP-element group 391: 	 branch_block_stmt_32/if_stmt_836_if_link/$entry
      -- CP-element group 391: 	 branch_block_stmt_32/if_stmt_836_else_link/$entry
      -- CP-element group 391: 	 branch_block_stmt_32/merge_stmt_819_PhiAck/$exit
      -- CP-element group 391: 	 branch_block_stmt_32/merge_stmt_819_PhiAck/$entry
      -- CP-element group 391: 	 branch_block_stmt_32/merge_stmt_819_PhiAck/dummy
      -- 
    branch_req_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(391), ack => if_stmt_836_branch_req_0); -- 
    convTranspose_CP_39_elements(391) <= OrReduce(convTranspose_CP_39_elements(188) & convTranspose_CP_39_elements(101));
    -- CP-element group 392:  transition  output  delay-element  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	193 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	396 
    -- CP-element group 392:  members (5) 
      -- CP-element group 392: 	 branch_block_stmt_32/bbx_xnph481_forx_xbody266_PhiReq/$exit
      -- CP-element group 392: 	 branch_block_stmt_32/bbx_xnph481_forx_xbody266_PhiReq/phi_stmt_880/$exit
      -- CP-element group 392: 	 branch_block_stmt_32/bbx_xnph481_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_req
      -- CP-element group 392: 	 branch_block_stmt_32/bbx_xnph481_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_sources/type_cast_886_konst_delay_trans
      -- CP-element group 392: 	 branch_block_stmt_32/bbx_xnph481_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_sources/$exit
      -- 
    phi_stmt_880_req_3128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_880_req_3128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(392), ack => phi_stmt_880_req_1); -- 
    -- Element group convTranspose_CP_39_elements(392) is a control-delay.
    cp_element_392_delay: control_delay_element  generic map(name => " 392_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(193), ack => convTranspose_CP_39_elements(392), clk => clk, reset =>reset);
    -- CP-element group 393:  transition  input  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	202 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	395 
    -- CP-element group 393:  members (2) 
      -- CP-element group 393: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_sources/type_cast_883/SplitProtocol/Sample/$exit
      -- CP-element group 393: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_sources/type_cast_883/SplitProtocol/Sample/ra
      -- 
    ra_3148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_883_inst_ack_0, ack => convTranspose_CP_39_elements(393)); -- 
    -- CP-element group 394:  transition  input  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	202 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	395 
    -- CP-element group 394:  members (2) 
      -- CP-element group 394: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_sources/type_cast_883/SplitProtocol/Update/ca
      -- CP-element group 394: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_sources/type_cast_883/SplitProtocol/Update/$exit
      -- 
    ca_3153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_883_inst_ack_1, ack => convTranspose_CP_39_elements(394)); -- 
    -- CP-element group 395:  join  transition  output  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	393 
    -- CP-element group 395: 	394 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	396 
    -- CP-element group 395:  members (6) 
      -- CP-element group 395: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_sources/type_cast_883/SplitProtocol/$exit
      -- CP-element group 395: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_sources/type_cast_883/$exit
      -- CP-element group 395: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_sources/$exit
      -- CP-element group 395: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_880/$exit
      -- CP-element group 395: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/$exit
      -- CP-element group 395: 	 branch_block_stmt_32/forx_xbody266_forx_xbody266_PhiReq/phi_stmt_880/phi_stmt_880_req
      -- 
    phi_stmt_880_req_3154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_880_req_3154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(395), ack => phi_stmt_880_req_0); -- 
    convTranspose_cp_element_group_395: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_395"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(393) & convTranspose_CP_39_elements(394);
      gj_convTranspose_cp_element_group_395 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(395), clk => clk, reset => reset); --
    end block;
    -- CP-element group 396:  merge  transition  place  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	392 
    -- CP-element group 396: 	395 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	397 
    -- CP-element group 396:  members (2) 
      -- CP-element group 396: 	 branch_block_stmt_32/merge_stmt_879_PhiReqMerge
      -- CP-element group 396: 	 branch_block_stmt_32/merge_stmt_879_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(396) <= OrReduce(convTranspose_CP_39_elements(392) & convTranspose_CP_39_elements(395));
    -- CP-element group 397:  fork  transition  place  input  output  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	396 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	194 
    -- CP-element group 397: 	195 
    -- CP-element group 397: 	197 
    -- CP-element group 397: 	199 
    -- CP-element group 397:  members (29) 
      -- CP-element group 397: 	 branch_block_stmt_32/merge_stmt_879__exit__
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910__entry__
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/$entry
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/addr_of_893_update_start_
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_index_resized_1
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_index_scaled_1
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_index_computed_1
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_index_resize_1/$entry
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_index_resize_1/$exit
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_index_resize_1/index_resize_req
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_index_resize_1/index_resize_ack
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_index_scale_1/$entry
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_index_scale_1/$exit
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_index_scale_1/scale_rename_req
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_index_scale_1/scale_rename_ack
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_final_index_sum_regn_update_start
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_final_index_sum_regn_Sample/$entry
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_final_index_sum_regn_Sample/req
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_final_index_sum_regn_Update/$entry
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/array_obj_ref_892_final_index_sum_regn_Update/req
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/addr_of_893_complete/$entry
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/addr_of_893_complete/req
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_update_start_
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Update/$entry
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Update/word_access_complete/$entry
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Update/word_access_complete/word_0/$entry
      -- CP-element group 397: 	 branch_block_stmt_32/assign_stmt_894_to_assign_stmt_910/ptr_deref_896_Update/word_access_complete/word_0/cr
      -- CP-element group 397: 	 branch_block_stmt_32/merge_stmt_879_PhiAck/phi_stmt_880_ack
      -- CP-element group 397: 	 branch_block_stmt_32/merge_stmt_879_PhiAck/$exit
      -- 
    phi_stmt_880_ack_3159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_880_ack_0, ack => convTranspose_CP_39_elements(397)); -- 
    req_1623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(397), ack => array_obj_ref_892_index_offset_req_0); -- 
    req_1628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(397), ack => array_obj_ref_892_index_offset_req_1); -- 
    req_1643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(397), ack => addr_of_893_final_reg_req_1); -- 
    cr_1693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(397), ack => ptr_deref_896_store_0_req_1); -- 
    -- CP-element group 398:  merge  fork  transition  place  output  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	191 
    -- CP-element group 398: 	201 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	203 
    -- CP-element group 398: 	204 
    -- CP-element group 398: 	206 
    -- CP-element group 398: 	207 
    -- CP-element group 398: 	233 
    -- CP-element group 398: 	259 
    -- CP-element group 398: 	285 
    -- CP-element group 398: 	311 
    -- CP-element group 398: 	313 
    -- CP-element group 398: 	315 
    -- CP-element group 398: 	317 
    -- CP-element group 398:  members (40) 
      -- CP-element group 398: 	 branch_block_stmt_32/merge_stmt_919__exit__
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097__entry__
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1008_sample_start_
      -- CP-element group 398: 	 branch_block_stmt_32/merge_stmt_919_PhiReqMerge
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1008_Sample/$entry
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block2_start_1008_Sample/req
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1047_Sample/req
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1047_Sample/$entry
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block3_start_1047_sample_start_
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/$entry
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/call_stmt_922_sample_start_
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/call_stmt_922_update_start_
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/call_stmt_922_Sample/$entry
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/call_stmt_922_Sample/crr
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/call_stmt_922_Update/$entry
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/call_stmt_922_Update/ccr
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/type_cast_927_update_start_
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/type_cast_927_Update/$entry
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/type_cast_927_Update/cr
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_929_sample_start_
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_929_Sample/$entry
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block0_start_929_Sample/req
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_969_sample_start_
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_969_Sample/$entry
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/WPIPE_Block1_start_969_Sample/req
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block0_done_1087_sample_start_
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block0_done_1087_Sample/$entry
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block0_done_1087_Sample/rr
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block1_done_1090_sample_start_
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block1_done_1090_Sample/$entry
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block1_done_1090_Sample/rr
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block2_done_1093_sample_start_
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block2_done_1093_Sample/$entry
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block2_done_1093_Sample/rr
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block3_done_1096_sample_start_
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block3_done_1096_Sample/$entry
      -- CP-element group 398: 	 branch_block_stmt_32/call_stmt_922_to_assign_stmt_1097/RPIPE_Block3_done_1096_Sample/rr
      -- CP-element group 398: 	 branch_block_stmt_32/merge_stmt_919_PhiAck/dummy
      -- CP-element group 398: 	 branch_block_stmt_32/merge_stmt_919_PhiAck/$exit
      -- CP-element group 398: 	 branch_block_stmt_32/merge_stmt_919_PhiAck/$entry
      -- 
    req_2116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(398), ack => WPIPE_Block2_start_1008_inst_req_0); -- 
    req_2298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(398), ack => WPIPE_Block3_start_1047_inst_req_0); -- 
    crr_1724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(398), ack => call_stmt_922_call_req_0); -- 
    ccr_1729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(398), ack => call_stmt_922_call_req_1); -- 
    cr_1743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(398), ack => type_cast_927_inst_req_1); -- 
    req_1752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(398), ack => WPIPE_Block0_start_929_inst_req_0); -- 
    req_1934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(398), ack => WPIPE_Block1_start_969_inst_req_0); -- 
    rr_2480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(398), ack => RPIPE_Block0_done_1087_inst_req_0); -- 
    rr_2494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(398), ack => RPIPE_Block1_done_1090_inst_req_0); -- 
    rr_2508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(398), ack => RPIPE_Block2_done_1093_inst_req_0); -- 
    rr_2522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(398), ack => RPIPE_Block3_done_1096_inst_req_0); -- 
    convTranspose_CP_39_elements(398) <= OrReduce(convTranspose_CP_39_elements(191) & convTranspose_CP_39_elements(201));
    -- CP-element group 399:  transition  output  delay-element  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	329 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	403 
    -- CP-element group 399:  members (5) 
      -- CP-element group 399: 	 branch_block_stmt_32/bbx_xnph_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_req
      -- CP-element group 399: 	 branch_block_stmt_32/bbx_xnph_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_sources/type_cast_1165_konst_delay_trans
      -- CP-element group 399: 	 branch_block_stmt_32/bbx_xnph_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_sources/$exit
      -- CP-element group 399: 	 branch_block_stmt_32/bbx_xnph_forx_xbody402_PhiReq/phi_stmt_1159/$exit
      -- CP-element group 399: 	 branch_block_stmt_32/bbx_xnph_forx_xbody402_PhiReq/$exit
      -- 
    phi_stmt_1159_req_3205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1159_req_3205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(399), ack => phi_stmt_1159_req_1); -- 
    -- Element group convTranspose_CP_39_elements(399) is a control-delay.
    cp_element_399_delay: control_delay_element  generic map(name => " 399_delay", delay_value => 1)  port map(req => convTranspose_CP_39_elements(329), ack => convTranspose_CP_39_elements(399), clk => clk, reset =>reset);
    -- CP-element group 400:  transition  input  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	377 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	402 
    -- CP-element group 400:  members (2) 
      -- CP-element group 400: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_sources/type_cast_1162/SplitProtocol/Sample/ra
      -- CP-element group 400: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_sources/type_cast_1162/SplitProtocol/Sample/$exit
      -- 
    ra_3225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1162_inst_ack_0, ack => convTranspose_CP_39_elements(400)); -- 
    -- CP-element group 401:  transition  input  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	377 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	402 
    -- CP-element group 401:  members (2) 
      -- CP-element group 401: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_sources/type_cast_1162/SplitProtocol/Update/$exit
      -- CP-element group 401: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_sources/type_cast_1162/SplitProtocol/Update/ca
      -- 
    ca_3230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1162_inst_ack_1, ack => convTranspose_CP_39_elements(401)); -- 
    -- CP-element group 402:  join  transition  output  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	400 
    -- CP-element group 402: 	401 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	403 
    -- CP-element group 402:  members (6) 
      -- CP-element group 402: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_sources/type_cast_1162/$exit
      -- CP-element group 402: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_sources/type_cast_1162/SplitProtocol/$exit
      -- CP-element group 402: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_req
      -- CP-element group 402: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/phi_stmt_1159/phi_stmt_1159_sources/$exit
      -- CP-element group 402: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/phi_stmt_1159/$exit
      -- CP-element group 402: 	 branch_block_stmt_32/forx_xbody402_forx_xbody402_PhiReq/$exit
      -- 
    phi_stmt_1159_req_3231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1159_req_3231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(402), ack => phi_stmt_1159_req_0); -- 
    convTranspose_cp_element_group_402: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTranspose_cp_element_group_402"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_39_elements(400) & convTranspose_CP_39_elements(401);
      gj_convTranspose_cp_element_group_402 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_39_elements(402), clk => clk, reset => reset); --
    end block;
    -- CP-element group 403:  merge  transition  place  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	399 
    -- CP-element group 403: 	402 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	404 
    -- CP-element group 403:  members (2) 
      -- CP-element group 403: 	 branch_block_stmt_32/merge_stmt_1158_PhiReqMerge
      -- CP-element group 403: 	 branch_block_stmt_32/merge_stmt_1158_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(403) <= OrReduce(convTranspose_CP_39_elements(399) & convTranspose_CP_39_elements(402));
    -- CP-element group 404:  fork  transition  place  input  output  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	403 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	330 
    -- CP-element group 404: 	331 
    -- CP-element group 404: 	333 
    -- CP-element group 404: 	335 
    -- CP-element group 404: 	337 
    -- CP-element group 404: 	339 
    -- CP-element group 404: 	341 
    -- CP-element group 404: 	343 
    -- CP-element group 404: 	345 
    -- CP-element group 404: 	347 
    -- CP-element group 404: 	349 
    -- CP-element group 404: 	351 
    -- CP-element group 404:  members (53) 
      -- CP-element group 404: 	 branch_block_stmt_32/merge_stmt_1158__exit__
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286__entry__
      -- CP-element group 404: 	 branch_block_stmt_32/merge_stmt_1158_PhiAck/$exit
      -- CP-element group 404: 	 branch_block_stmt_32/merge_stmt_1158_PhiAck/phi_stmt_1159_ack
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/addr_of_1172_update_start_
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_index_resized_1
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_index_scaled_1
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_index_computed_1
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_index_resize_1/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_index_resize_1/$exit
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_index_resize_1/index_resize_req
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_index_resize_1/index_resize_ack
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_index_scale_1/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_index_scale_1/$exit
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_index_scale_1/scale_rename_req
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_index_scale_1/scale_rename_ack
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_final_index_sum_regn_update_start
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_final_index_sum_regn_Sample/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_final_index_sum_regn_Sample/req
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_final_index_sum_regn_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/array_obj_ref_1171_final_index_sum_regn_Update/req
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/addr_of_1172_complete/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/addr_of_1172_complete/req
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_update_start_
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Update/word_access_complete/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Update/word_access_complete/word_0/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/ptr_deref_1176_Update/word_access_complete/word_0/cr
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1180_update_start_
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1180_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1180_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1190_update_start_
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1190_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1190_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1200_update_start_
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1200_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1200_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1210_update_start_
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1210_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1210_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1220_update_start_
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1220_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1220_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1230_update_start_
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1230_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1230_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1240_update_start_
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1240_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1240_Update/cr
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1250_update_start_
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1250_Update/$entry
      -- CP-element group 404: 	 branch_block_stmt_32/assign_stmt_1173_to_assign_stmt_1286/type_cast_1250_Update/cr
      -- 
    phi_stmt_1159_ack_3236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1159_ack_0, ack => convTranspose_CP_39_elements(404)); -- 
    req_2637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => array_obj_ref_1171_index_offset_req_0); -- 
    req_2642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => array_obj_ref_1171_index_offset_req_1); -- 
    req_2657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => addr_of_1172_final_reg_req_1); -- 
    cr_2702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => ptr_deref_1176_load_0_req_1); -- 
    cr_2721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_1180_inst_req_1); -- 
    cr_2735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_1190_inst_req_1); -- 
    cr_2749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_1200_inst_req_1); -- 
    cr_2763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_1210_inst_req_1); -- 
    cr_2777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_1220_inst_req_1); -- 
    cr_2791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_1230_inst_req_1); -- 
    cr_2805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_1240_inst_req_1); -- 
    cr_2819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_39_elements(404), ack => type_cast_1250_inst_req_1); -- 
    -- CP-element group 405:  merge  transition  place  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	327 
    -- CP-element group 405: 	376 
    -- CP-element group 405: successors 
    -- CP-element group 405:  members (16) 
      -- CP-element group 405: 	 $exit
      -- CP-element group 405: 	 branch_block_stmt_32/$exit
      -- CP-element group 405: 	 branch_block_stmt_32/branch_block_stmt_32__exit__
      -- CP-element group 405: 	 branch_block_stmt_32/merge_stmt_1295__exit__
      -- CP-element group 405: 	 branch_block_stmt_32/return__
      -- CP-element group 405: 	 branch_block_stmt_32/merge_stmt_1297__exit__
      -- CP-element group 405: 	 branch_block_stmt_32/merge_stmt_1295_PhiReqMerge
      -- CP-element group 405: 	 branch_block_stmt_32/merge_stmt_1297_PhiReqMerge
      -- CP-element group 405: 	 branch_block_stmt_32/merge_stmt_1297_PhiAck/dummy
      -- CP-element group 405: 	 branch_block_stmt_32/merge_stmt_1297_PhiAck/$exit
      -- CP-element group 405: 	 branch_block_stmt_32/merge_stmt_1297_PhiAck/$entry
      -- CP-element group 405: 	 branch_block_stmt_32/return___PhiReq/$exit
      -- CP-element group 405: 	 branch_block_stmt_32/return___PhiReq/$entry
      -- CP-element group 405: 	 branch_block_stmt_32/merge_stmt_1295_PhiAck/dummy
      -- CP-element group 405: 	 branch_block_stmt_32/merge_stmt_1295_PhiAck/$exit
      -- CP-element group 405: 	 branch_block_stmt_32/merge_stmt_1295_PhiAck/$entry
      -- 
    convTranspose_CP_39_elements(405) <= OrReduce(convTranspose_CP_39_elements(327) & convTranspose_CP_39_elements(376));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar499_891_resized : std_logic_vector(13 downto 0);
    signal R_indvar499_891_scaled : std_logic_vector(13 downto 0);
    signal R_indvar513_659_resized : std_logic_vector(10 downto 0);
    signal R_indvar513_659_scaled : std_logic_vector(10 downto 0);
    signal R_indvar529_452_resized : std_logic_vector(13 downto 0);
    signal R_indvar529_452_scaled : std_logic_vector(13 downto 0);
    signal R_indvar_1170_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1170_scaled : std_logic_vector(13 downto 0);
    signal add108_305 : std_logic_vector(31 downto 0);
    signal add117_330 : std_logic_vector(31 downto 0);
    signal add126_355 : std_logic_vector(31 downto 0);
    signal add12_82 : std_logic_vector(31 downto 0);
    signal add135_380 : std_logic_vector(31 downto 0);
    signal add150_480 : std_logic_vector(63 downto 0);
    signal add156_498 : std_logic_vector(63 downto 0);
    signal add162_516 : std_logic_vector(63 downto 0);
    signal add168_534 : std_logic_vector(63 downto 0);
    signal add174_552 : std_logic_vector(63 downto 0);
    signal add180_570 : std_logic_vector(63 downto 0);
    signal add186_588 : std_logic_vector(63 downto 0);
    signal add206_687 : std_logic_vector(63 downto 0);
    signal add212_705 : std_logic_vector(63 downto 0);
    signal add218_723 : std_logic_vector(63 downto 0);
    signal add21_107 : std_logic_vector(31 downto 0);
    signal add224_741 : std_logic_vector(63 downto 0);
    signal add230_759 : std_logic_vector(63 downto 0);
    signal add236_777 : std_logic_vector(63 downto 0);
    signal add242_795 : std_logic_vector(63 downto 0);
    signal add30_132 : std_logic_vector(31 downto 0);
    signal add39_157 : std_logic_vector(31 downto 0);
    signal add48_182 : std_logic_vector(31 downto 0);
    signal add57_207 : std_logic_vector(31 downto 0);
    signal add74_235 : std_logic_vector(31 downto 0);
    signal add79_240 : std_logic_vector(31 downto 0);
    signal add99_280 : std_logic_vector(31 downto 0);
    signal add_57 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1171_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1171_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1171_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1171_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1171_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1171_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_453_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_453_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_453_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_453_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_453_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_453_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_660_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_660_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_660_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_660_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_660_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_660_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_892_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_892_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_892_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_892_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_892_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_892_root_address : std_logic_vector(13 downto 0);
    signal arrayidx246_662 : std_logic_vector(31 downto 0);
    signal arrayidx269_894 : std_logic_vector(31 downto 0);
    signal arrayidx407_1173 : std_logic_vector(31 downto 0);
    signal arrayidx_455 : std_logic_vector(31 downto 0);
    signal call101_283 : std_logic_vector(7 downto 0);
    signal call106_296 : std_logic_vector(7 downto 0);
    signal call10_73 : std_logic_vector(7 downto 0);
    signal call110_308 : std_logic_vector(7 downto 0);
    signal call115_321 : std_logic_vector(7 downto 0);
    signal call119_333 : std_logic_vector(7 downto 0);
    signal call124_346 : std_logic_vector(7 downto 0);
    signal call128_358 : std_logic_vector(7 downto 0);
    signal call133_371 : std_logic_vector(7 downto 0);
    signal call143_458 : std_logic_vector(7 downto 0);
    signal call147_471 : std_logic_vector(7 downto 0);
    signal call14_85 : std_logic_vector(7 downto 0);
    signal call153_489 : std_logic_vector(7 downto 0);
    signal call159_507 : std_logic_vector(7 downto 0);
    signal call165_525 : std_logic_vector(7 downto 0);
    signal call171_543 : std_logic_vector(7 downto 0);
    signal call177_561 : std_logic_vector(7 downto 0);
    signal call183_579 : std_logic_vector(7 downto 0);
    signal call199_665 : std_logic_vector(7 downto 0);
    signal call19_98 : std_logic_vector(7 downto 0);
    signal call203_678 : std_logic_vector(7 downto 0);
    signal call209_696 : std_logic_vector(7 downto 0);
    signal call215_714 : std_logic_vector(7 downto 0);
    signal call221_732 : std_logic_vector(7 downto 0);
    signal call227_750 : std_logic_vector(7 downto 0);
    signal call233_768 : std_logic_vector(7 downto 0);
    signal call239_786 : std_logic_vector(7 downto 0);
    signal call23_110 : std_logic_vector(7 downto 0);
    signal call275_922 : std_logic_vector(63 downto 0);
    signal call28_123 : std_logic_vector(7 downto 0);
    signal call2_48 : std_logic_vector(7 downto 0);
    signal call32_135 : std_logic_vector(7 downto 0);
    signal call378_1088 : std_logic_vector(31 downto 0);
    signal call37_148 : std_logic_vector(7 downto 0);
    signal call381_1091 : std_logic_vector(31 downto 0);
    signal call384_1094 : std_logic_vector(31 downto 0);
    signal call387_1097 : std_logic_vector(31 downto 0);
    signal call390_1100 : std_logic_vector(63 downto 0);
    signal call41_160 : std_logic_vector(7 downto 0);
    signal call46_173 : std_logic_vector(7 downto 0);
    signal call50_185 : std_logic_vector(7 downto 0);
    signal call55_198 : std_logic_vector(7 downto 0);
    signal call5_60 : std_logic_vector(7 downto 0);
    signal call92_258 : std_logic_vector(7 downto 0);
    signal call97_271 : std_logic_vector(7 downto 0);
    signal call_35 : std_logic_vector(7 downto 0);
    signal cmp194483_402 : std_logic_vector(0 downto 0);
    signal cmp264479_835 : std_logic_vector(0 downto 0);
    signal cmp487_387 : std_logic_vector(0 downto 0);
    signal conv104_287 : std_logic_vector(31 downto 0);
    signal conv107_300 : std_logic_vector(31 downto 0);
    signal conv113_312 : std_logic_vector(31 downto 0);
    signal conv116_325 : std_logic_vector(31 downto 0);
    signal conv11_77 : std_logic_vector(31 downto 0);
    signal conv122_337 : std_logic_vector(31 downto 0);
    signal conv125_350 : std_logic_vector(31 downto 0);
    signal conv131_362 : std_logic_vector(31 downto 0);
    signal conv134_375 : std_logic_vector(31 downto 0);
    signal conv144_462 : std_logic_vector(63 downto 0);
    signal conv149_475 : std_logic_vector(63 downto 0);
    signal conv155_493 : std_logic_vector(63 downto 0);
    signal conv161_511 : std_logic_vector(63 downto 0);
    signal conv167_529 : std_logic_vector(63 downto 0);
    signal conv173_547 : std_logic_vector(63 downto 0);
    signal conv179_565 : std_logic_vector(63 downto 0);
    signal conv17_89 : std_logic_vector(31 downto 0);
    signal conv185_583 : std_logic_vector(63 downto 0);
    signal conv1_39 : std_logic_vector(31 downto 0);
    signal conv200_669 : std_logic_vector(63 downto 0);
    signal conv205_682 : std_logic_vector(63 downto 0);
    signal conv20_102 : std_logic_vector(31 downto 0);
    signal conv211_700 : std_logic_vector(63 downto 0);
    signal conv217_718 : std_logic_vector(63 downto 0);
    signal conv223_736 : std_logic_vector(63 downto 0);
    signal conv229_754 : std_logic_vector(63 downto 0);
    signal conv235_772 : std_logic_vector(63 downto 0);
    signal conv241_790 : std_logic_vector(63 downto 0);
    signal conv26_114 : std_logic_vector(31 downto 0);
    signal conv276_928 : std_logic_vector(63 downto 0);
    signal conv29_127 : std_logic_vector(31 downto 0);
    signal conv35_139 : std_logic_vector(31 downto 0);
    signal conv38_152 : std_logic_vector(31 downto 0);
    signal conv391_1105 : std_logic_vector(63 downto 0);
    signal conv3_52 : std_logic_vector(31 downto 0);
    signal conv411_1181 : std_logic_vector(7 downto 0);
    signal conv417_1191 : std_logic_vector(7 downto 0);
    signal conv423_1201 : std_logic_vector(7 downto 0);
    signal conv429_1211 : std_logic_vector(7 downto 0);
    signal conv435_1221 : std_logic_vector(7 downto 0);
    signal conv441_1231 : std_logic_vector(7 downto 0);
    signal conv447_1241 : std_logic_vector(7 downto 0);
    signal conv44_164 : std_logic_vector(31 downto 0);
    signal conv453_1251 : std_logic_vector(7 downto 0);
    signal conv47_177 : std_logic_vector(31 downto 0);
    signal conv53_189 : std_logic_vector(31 downto 0);
    signal conv56_202 : std_logic_vector(31 downto 0);
    signal conv8_64 : std_logic_vector(31 downto 0);
    signal conv95_262 : std_logic_vector(31 downto 0);
    signal conv98_275 : std_logic_vector(31 downto 0);
    signal exitcond1_1286 : std_logic_vector(0 downto 0);
    signal exitcond2_810 : std_logic_vector(0 downto 0);
    signal exitcond3_603 : std_logic_vector(0 downto 0);
    signal exitcond_910 : std_logic_vector(0 downto 0);
    signal iNsTr_14_229 : std_logic_vector(31 downto 0);
    signal iNsTr_172_1143 : std_logic_vector(63 downto 0);
    signal iNsTr_26_425 : std_logic_vector(63 downto 0);
    signal iNsTr_39_632 : std_logic_vector(63 downto 0);
    signal iNsTr_53_864 : std_logic_vector(63 downto 0);
    signal indvar499_880 : std_logic_vector(63 downto 0);
    signal indvar513_648 : std_logic_vector(63 downto 0);
    signal indvar529_441 : std_logic_vector(63 downto 0);
    signal indvar_1159 : std_logic_vector(63 downto 0);
    signal indvarx_xnext500_905 : std_logic_vector(63 downto 0);
    signal indvarx_xnext514_805 : std_logic_vector(63 downto 0);
    signal indvarx_xnext530_598 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1281 : std_logic_vector(63 downto 0);
    signal mul256_824 : std_logic_vector(31 downto 0);
    signal mul259_829 : std_logic_vector(31 downto 0);
    signal mul66_217 : std_logic_vector(31 downto 0);
    signal mul85_245 : std_logic_vector(31 downto 0);
    signal mul88_250 : std_logic_vector(31 downto 0);
    signal mul91_255 : std_logic_vector(31 downto 0);
    signal mul_212 : std_logic_vector(31 downto 0);
    signal ptr_deref_1176_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1176_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1176_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1176_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1176_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_590_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_590_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_590_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_590_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_590_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_590_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_797_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_797_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_797_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_797_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_797_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_797_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_896_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_896_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_896_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_896_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_896_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_896_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl105_293 : std_logic_vector(31 downto 0);
    signal shl114_318 : std_logic_vector(31 downto 0);
    signal shl123_343 : std_logic_vector(31 downto 0);
    signal shl132_368 : std_logic_vector(31 downto 0);
    signal shl146_468 : std_logic_vector(63 downto 0);
    signal shl152_486 : std_logic_vector(63 downto 0);
    signal shl158_504 : std_logic_vector(63 downto 0);
    signal shl164_522 : std_logic_vector(63 downto 0);
    signal shl170_540 : std_logic_vector(63 downto 0);
    signal shl176_558 : std_logic_vector(63 downto 0);
    signal shl182_576 : std_logic_vector(63 downto 0);
    signal shl18_95 : std_logic_vector(31 downto 0);
    signal shl202_675 : std_logic_vector(63 downto 0);
    signal shl208_693 : std_logic_vector(63 downto 0);
    signal shl214_711 : std_logic_vector(63 downto 0);
    signal shl220_729 : std_logic_vector(63 downto 0);
    signal shl226_747 : std_logic_vector(63 downto 0);
    signal shl232_765 : std_logic_vector(63 downto 0);
    signal shl238_783 : std_logic_vector(63 downto 0);
    signal shl27_120 : std_logic_vector(31 downto 0);
    signal shl36_145 : std_logic_vector(31 downto 0);
    signal shl45_170 : std_logic_vector(31 downto 0);
    signal shl54_195 : std_logic_vector(31 downto 0);
    signal shl96_268 : std_logic_vector(31 downto 0);
    signal shl9_70 : std_logic_vector(31 downto 0);
    signal shl_45 : std_logic_vector(31 downto 0);
    signal shr414_1187 : std_logic_vector(63 downto 0);
    signal shr420_1197 : std_logic_vector(63 downto 0);
    signal shr426_1207 : std_logic_vector(63 downto 0);
    signal shr432_1217 : std_logic_vector(63 downto 0);
    signal shr438_1227 : std_logic_vector(63 downto 0);
    signal shr444_1237 : std_logic_vector(63 downto 0);
    signal shr450_1247 : std_logic_vector(63 downto 0);
    signal shr_223 : std_logic_vector(31 downto 0);
    signal sub_1110 : std_logic_vector(63 downto 0);
    signal tmp408_1177 : std_logic_vector(63 downto 0);
    signal tmp494_1127 : std_logic_vector(31 downto 0);
    signal tmp494x_xop_1139 : std_logic_vector(31 downto 0);
    signal tmp495_1133 : std_logic_vector(0 downto 0);
    signal tmp498_1156 : std_logic_vector(63 downto 0);
    signal tmp506_848 : std_logic_vector(31 downto 0);
    signal tmp506x_xop_860 : std_logic_vector(31 downto 0);
    signal tmp507_854 : std_logic_vector(0 downto 0);
    signal tmp511_877 : std_logic_vector(63 downto 0);
    signal tmp522_616 : std_logic_vector(31 downto 0);
    signal tmp522x_xop_628 : std_logic_vector(31 downto 0);
    signal tmp523_622 : std_logic_vector(0 downto 0);
    signal tmp527_645 : std_logic_vector(63 downto 0);
    signal tmp536x_xop_421 : std_logic_vector(31 downto 0);
    signal tmp537_415 : std_logic_vector(0 downto 0);
    signal tmp541_438 : std_logic_vector(63 downto 0);
    signal type_cast_1103_wire : std_logic_vector(63 downto 0);
    signal type_cast_1125_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1131_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1137_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1147_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1154_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1162_wire : std_logic_vector(63 downto 0);
    signal type_cast_1165_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1185_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_118_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1195_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1205_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1215_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1225_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1235_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1245_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1279_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_143_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_168_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_193_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_221_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_227_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_233_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_266_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_291_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_316_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_341_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_366_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_384_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_400_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_413_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_419_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_429_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_436_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_43_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_445_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_447_wire : std_logic_vector(63 downto 0);
    signal type_cast_466_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_484_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_502_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_520_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_538_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_556_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_574_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_596_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_614_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_620_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_626_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_636_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_643_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_651_wire : std_logic_vector(63 downto 0);
    signal type_cast_654_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_673_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_68_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_691_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_709_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_727_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_745_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_763_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_781_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_803_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_833_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_846_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_852_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_858_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_868_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_875_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_883_wire : std_logic_vector(63 downto 0);
    signal type_cast_886_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_898_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_903_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_926_wire : std_logic_vector(63 downto 0);
    signal type_cast_93_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_958_wire_constant : std_logic_vector(31 downto 0);
    signal xx_xop543_870 : std_logic_vector(63 downto 0);
    signal xx_xop544_638 : std_logic_vector(63 downto 0);
    signal xx_xop545_431 : std_logic_vector(63 downto 0);
    signal xx_xop_1149 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1171_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1171_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1171_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1171_resized_base_address <= "00000000000000";
    array_obj_ref_453_constant_part_of_offset <= "00000000000000";
    array_obj_ref_453_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_453_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_453_resized_base_address <= "00000000000000";
    array_obj_ref_660_constant_part_of_offset <= "00000100010";
    array_obj_ref_660_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_660_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_660_resized_base_address <= "00000000000";
    array_obj_ref_892_constant_part_of_offset <= "00000000000000";
    array_obj_ref_892_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_892_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_892_resized_base_address <= "00000000000000";
    ptr_deref_1176_word_offset_0 <= "00000000000000";
    ptr_deref_590_word_offset_0 <= "00000000000000";
    ptr_deref_797_word_offset_0 <= "00000000000";
    ptr_deref_896_word_offset_0 <= "00000000000000";
    type_cast_1125_wire_constant <= "00000000000000000000000000000010";
    type_cast_1131_wire_constant <= "00000000000000000000000000000001";
    type_cast_1137_wire_constant <= "11111111111111111111111111111111";
    type_cast_1147_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1154_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1165_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1185_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_118_wire_constant <= "00000000000000000000000000001000";
    type_cast_1195_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1205_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1215_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1225_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1235_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1245_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1279_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_143_wire_constant <= "00000000000000000000000000001000";
    type_cast_168_wire_constant <= "00000000000000000000000000001000";
    type_cast_193_wire_constant <= "00000000000000000000000000001000";
    type_cast_221_wire_constant <= "00000000000000000000000000000010";
    type_cast_227_wire_constant <= "00000000000000000000000000000001";
    type_cast_233_wire_constant <= "01111111111111111111111111111110";
    type_cast_266_wire_constant <= "00000000000000000000000000001000";
    type_cast_291_wire_constant <= "00000000000000000000000000001000";
    type_cast_316_wire_constant <= "00000000000000000000000000001000";
    type_cast_341_wire_constant <= "00000000000000000000000000001000";
    type_cast_366_wire_constant <= "00000000000000000000000000001000";
    type_cast_384_wire_constant <= "00000000000000000000000000000011";
    type_cast_400_wire_constant <= "00000000000000000000000000000011";
    type_cast_413_wire_constant <= "00000000000000000000000000000001";
    type_cast_419_wire_constant <= "11111111111111111111111111111111";
    type_cast_429_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_436_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_43_wire_constant <= "00000000000000000000000000001000";
    type_cast_445_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_466_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_484_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_502_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_520_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_538_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_556_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_574_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_596_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_614_wire_constant <= "00000000000000000000000000000010";
    type_cast_620_wire_constant <= "00000000000000000000000000000001";
    type_cast_626_wire_constant <= "11111111111111111111111111111111";
    type_cast_636_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_643_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_654_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_673_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_68_wire_constant <= "00000000000000000000000000001000";
    type_cast_691_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_709_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_727_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_745_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_763_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_781_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_803_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_833_wire_constant <= "00000000000000000000000000000011";
    type_cast_846_wire_constant <= "00000000000000000000000000000010";
    type_cast_852_wire_constant <= "00000000000000000000000000000001";
    type_cast_858_wire_constant <= "11111111111111111111111111111111";
    type_cast_868_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_875_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_886_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_898_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_903_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_93_wire_constant <= "00000000000000000000000000001000";
    type_cast_958_wire_constant <= "00000000000000000000000000000000";
    phi_stmt_1159: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1162_wire & type_cast_1165_wire_constant;
      req <= phi_stmt_1159_req_0 & phi_stmt_1159_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1159",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1159_ack_0,
          idata => idata,
          odata => indvar_1159,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1159
    phi_stmt_441: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_445_wire_constant & type_cast_447_wire;
      req <= phi_stmt_441_req_0 & phi_stmt_441_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_441",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_441_ack_0,
          idata => idata,
          odata => indvar529_441,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_441
    phi_stmt_648: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_651_wire & type_cast_654_wire_constant;
      req <= phi_stmt_648_req_0 & phi_stmt_648_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_648",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_648_ack_0,
          idata => idata,
          odata => indvar513_648,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_648
    phi_stmt_880: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_883_wire & type_cast_886_wire_constant;
      req <= phi_stmt_880_req_0 & phi_stmt_880_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_880",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_880_ack_0,
          idata => idata,
          odata => indvar499_880,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_880
    -- flow-through select operator MUX_1155_inst
    tmp498_1156 <= xx_xop_1149 when (tmp495_1133(0) /=  '0') else type_cast_1154_wire_constant;
    -- flow-through select operator MUX_437_inst
    tmp541_438 <= xx_xop545_431 when (tmp537_415(0) /=  '0') else type_cast_436_wire_constant;
    -- flow-through select operator MUX_644_inst
    tmp527_645 <= xx_xop544_638 when (tmp523_622(0) /=  '0') else type_cast_643_wire_constant;
    -- flow-through select operator MUX_876_inst
    tmp511_877 <= xx_xop543_870 when (tmp507_854(0) /=  '0') else type_cast_875_wire_constant;
    addr_of_1172_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1172_final_reg_req_0;
      addr_of_1172_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1172_final_reg_req_1;
      addr_of_1172_final_reg_ack_1<= rack(0);
      addr_of_1172_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1172_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1171_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx407_1173,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_454_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_454_final_reg_req_0;
      addr_of_454_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_454_final_reg_req_1;
      addr_of_454_final_reg_ack_1<= rack(0);
      addr_of_454_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_454_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_453_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_455,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_661_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_661_final_reg_req_0;
      addr_of_661_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_661_final_reg_req_1;
      addr_of_661_final_reg_ack_1<= rack(0);
      addr_of_661_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_661_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_660_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx246_662,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_893_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_893_final_reg_req_0;
      addr_of_893_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_893_final_reg_req_1;
      addr_of_893_final_reg_ack_1<= rack(0);
      addr_of_893_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_893_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_892_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx269_894,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_101_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_101_inst_req_0;
      type_cast_101_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_101_inst_req_1;
      type_cast_101_inst_ack_1<= rack(0);
      type_cast_101_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_101_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_98,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_102,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1104_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1104_inst_req_0;
      type_cast_1104_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1104_inst_req_1;
      type_cast_1104_inst_ack_1<= rack(0);
      type_cast_1104_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1104_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1103_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv391_1105,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_113_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_113_inst_req_0;
      type_cast_113_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_113_inst_req_1;
      type_cast_113_inst_ack_1<= rack(0);
      type_cast_113_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_113_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_110,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_114,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1142_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1142_inst_req_0;
      type_cast_1142_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1142_inst_req_1;
      type_cast_1142_inst_ack_1<= rack(0);
      type_cast_1142_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1142_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp494x_xop_1139,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_172_1143,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1162_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1162_inst_req_0;
      type_cast_1162_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1162_inst_req_1;
      type_cast_1162_inst_ack_1<= rack(0);
      type_cast_1162_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1162_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1281,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1162_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1180_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1180_inst_req_0;
      type_cast_1180_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1180_inst_req_1;
      type_cast_1180_inst_ack_1<= rack(0);
      type_cast_1180_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1180_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp408_1177,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv411_1181,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1190_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1190_inst_req_0;
      type_cast_1190_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1190_inst_req_1;
      type_cast_1190_inst_ack_1<= rack(0);
      type_cast_1190_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1190_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr414_1187,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv417_1191,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1200_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1200_inst_req_0;
      type_cast_1200_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1200_inst_req_1;
      type_cast_1200_inst_ack_1<= rack(0);
      type_cast_1200_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1200_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr420_1197,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv423_1201,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1210_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1210_inst_req_0;
      type_cast_1210_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1210_inst_req_1;
      type_cast_1210_inst_ack_1<= rack(0);
      type_cast_1210_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1210_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr426_1207,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv429_1211,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1220_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1220_inst_req_0;
      type_cast_1220_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1220_inst_req_1;
      type_cast_1220_inst_ack_1<= rack(0);
      type_cast_1220_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1220_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr432_1217,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv435_1221,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1230_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1230_inst_req_0;
      type_cast_1230_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1230_inst_req_1;
      type_cast_1230_inst_ack_1<= rack(0);
      type_cast_1230_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1230_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr438_1227,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv441_1231,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1240_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1240_inst_req_0;
      type_cast_1240_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1240_inst_req_1;
      type_cast_1240_inst_ack_1<= rack(0);
      type_cast_1240_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1240_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr444_1237,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv447_1241,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1250_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1250_inst_req_0;
      type_cast_1250_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1250_inst_req_1;
      type_cast_1250_inst_ack_1<= rack(0);
      type_cast_1250_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1250_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr450_1247,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv453_1251,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_126_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_126_inst_req_0;
      type_cast_126_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_126_inst_req_1;
      type_cast_126_inst_ack_1<= rack(0);
      type_cast_126_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_126_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_123,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_127,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_138_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_138_inst_req_0;
      type_cast_138_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_138_inst_req_1;
      type_cast_138_inst_ack_1<= rack(0);
      type_cast_138_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_138_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_135,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_139,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_151_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_151_inst_req_0;
      type_cast_151_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_151_inst_req_1;
      type_cast_151_inst_ack_1<= rack(0);
      type_cast_151_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_151_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_148,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_152,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_163_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_163_inst_req_0;
      type_cast_163_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_163_inst_req_1;
      type_cast_163_inst_ack_1<= rack(0);
      type_cast_163_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_163_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_160,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_164,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_176_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_176_inst_req_0;
      type_cast_176_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_176_inst_req_1;
      type_cast_176_inst_ack_1<= rack(0);
      type_cast_176_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_176_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_173,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_177,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_188_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_188_inst_req_0;
      type_cast_188_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_188_inst_req_1;
      type_cast_188_inst_ack_1<= rack(0);
      type_cast_188_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_188_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_185,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_189,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_201_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_201_inst_req_0;
      type_cast_201_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_201_inst_req_1;
      type_cast_201_inst_ack_1<= rack(0);
      type_cast_201_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_201_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_198,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_202,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_261_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_261_inst_req_0;
      type_cast_261_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_261_inst_req_1;
      type_cast_261_inst_ack_1<= rack(0);
      type_cast_261_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_261_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call92_258,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_262,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_274_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_274_inst_req_0;
      type_cast_274_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_274_inst_req_1;
      type_cast_274_inst_ack_1<= rack(0);
      type_cast_274_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_274_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_271,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_275,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_286_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_286_inst_req_0;
      type_cast_286_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_286_inst_req_1;
      type_cast_286_inst_ack_1<= rack(0);
      type_cast_286_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_286_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_283,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_287,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_299_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_299_inst_req_0;
      type_cast_299_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_299_inst_req_1;
      type_cast_299_inst_ack_1<= rack(0);
      type_cast_299_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_299_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call106_296,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_300,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_311_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_311_inst_req_0;
      type_cast_311_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_311_inst_req_1;
      type_cast_311_inst_ack_1<= rack(0);
      type_cast_311_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_311_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call110_308,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_312,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_324_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_324_inst_req_0;
      type_cast_324_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_324_inst_req_1;
      type_cast_324_inst_ack_1<= rack(0);
      type_cast_324_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_324_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_321,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_325,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_336_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_336_inst_req_0;
      type_cast_336_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_336_inst_req_1;
      type_cast_336_inst_ack_1<= rack(0);
      type_cast_336_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_336_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_333,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_337,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_349_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_349_inst_req_0;
      type_cast_349_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_349_inst_req_1;
      type_cast_349_inst_ack_1<= rack(0);
      type_cast_349_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_349_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call124_346,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_350,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_361_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_361_inst_req_0;
      type_cast_361_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_361_inst_req_1;
      type_cast_361_inst_ack_1<= rack(0);
      type_cast_361_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_361_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_358,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_362,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_374_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_374_inst_req_0;
      type_cast_374_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_374_inst_req_1;
      type_cast_374_inst_ack_1<= rack(0);
      type_cast_374_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_374_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_371,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_375,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_38_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_38_inst_req_0;
      type_cast_38_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_38_inst_req_1;
      type_cast_38_inst_ack_1<= rack(0);
      type_cast_38_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_38_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_35,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_39,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_424_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_424_inst_req_0;
      type_cast_424_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_424_inst_req_1;
      type_cast_424_inst_ack_1<= rack(0);
      type_cast_424_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_424_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp536x_xop_421,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_26_425,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_447_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_447_inst_req_0;
      type_cast_447_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_447_inst_req_1;
      type_cast_447_inst_ack_1<= rack(0);
      type_cast_447_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_447_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext530_598,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_447_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_461_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_461_inst_req_0;
      type_cast_461_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_461_inst_req_1;
      type_cast_461_inst_ack_1<= rack(0);
      type_cast_461_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_461_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call143_458,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv144_462,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_474_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_474_inst_req_0;
      type_cast_474_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_474_inst_req_1;
      type_cast_474_inst_ack_1<= rack(0);
      type_cast_474_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_474_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call147_471,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv149_475,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_492_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_492_inst_req_0;
      type_cast_492_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_492_inst_req_1;
      type_cast_492_inst_ack_1<= rack(0);
      type_cast_492_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_492_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call153_489,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv155_493,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_510_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_510_inst_req_0;
      type_cast_510_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_510_inst_req_1;
      type_cast_510_inst_ack_1<= rack(0);
      type_cast_510_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_510_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call159_507,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv161_511,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_51_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_51_inst_req_0;
      type_cast_51_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_51_inst_req_1;
      type_cast_51_inst_ack_1<= rack(0);
      type_cast_51_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_51_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_48,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_52,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_528_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_528_inst_req_0;
      type_cast_528_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_528_inst_req_1;
      type_cast_528_inst_ack_1<= rack(0);
      type_cast_528_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_528_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call165_525,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv167_529,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_546_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_546_inst_req_0;
      type_cast_546_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_546_inst_req_1;
      type_cast_546_inst_ack_1<= rack(0);
      type_cast_546_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_546_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call171_543,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv173_547,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_564_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_564_inst_req_0;
      type_cast_564_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_564_inst_req_1;
      type_cast_564_inst_ack_1<= rack(0);
      type_cast_564_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_564_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call177_561,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv179_565,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_582_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_582_inst_req_0;
      type_cast_582_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_582_inst_req_1;
      type_cast_582_inst_ack_1<= rack(0);
      type_cast_582_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_582_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call183_579,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv185_583,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_631_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_631_inst_req_0;
      type_cast_631_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_631_inst_req_1;
      type_cast_631_inst_ack_1<= rack(0);
      type_cast_631_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_631_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp522x_xop_628,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_39_632,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_63_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_63_inst_req_0;
      type_cast_63_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_63_inst_req_1;
      type_cast_63_inst_ack_1<= rack(0);
      type_cast_63_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_63_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_60,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_64,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_651_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_651_inst_req_0;
      type_cast_651_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_651_inst_req_1;
      type_cast_651_inst_ack_1<= rack(0);
      type_cast_651_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_651_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext514_805,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_651_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_668_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_668_inst_req_0;
      type_cast_668_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_668_inst_req_1;
      type_cast_668_inst_ack_1<= rack(0);
      type_cast_668_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_668_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call199_665,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_669,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_681_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_681_inst_req_0;
      type_cast_681_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_681_inst_req_1;
      type_cast_681_inst_ack_1<= rack(0);
      type_cast_681_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_681_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call203_678,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv205_682,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_699_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_699_inst_req_0;
      type_cast_699_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_699_inst_req_1;
      type_cast_699_inst_ack_1<= rack(0);
      type_cast_699_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_699_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call209_696,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv211_700,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_717_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_717_inst_req_0;
      type_cast_717_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_717_inst_req_1;
      type_cast_717_inst_ack_1<= rack(0);
      type_cast_717_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_717_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call215_714,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv217_718,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_735_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_735_inst_req_0;
      type_cast_735_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_735_inst_req_1;
      type_cast_735_inst_ack_1<= rack(0);
      type_cast_735_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_735_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call221_732,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv223_736,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_753_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_753_inst_req_0;
      type_cast_753_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_753_inst_req_1;
      type_cast_753_inst_ack_1<= rack(0);
      type_cast_753_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_753_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call227_750,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv229_754,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_76_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_76_inst_req_0;
      type_cast_76_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_76_inst_req_1;
      type_cast_76_inst_ack_1<= rack(0);
      type_cast_76_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_76_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_73,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_77,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_771_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_771_inst_req_0;
      type_cast_771_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_771_inst_req_1;
      type_cast_771_inst_ack_1<= rack(0);
      type_cast_771_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_771_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call233_768,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv235_772,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_789_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_789_inst_req_0;
      type_cast_789_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_789_inst_req_1;
      type_cast_789_inst_ack_1<= rack(0);
      type_cast_789_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_789_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call239_786,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_790,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_863_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_863_inst_req_0;
      type_cast_863_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_863_inst_req_1;
      type_cast_863_inst_ack_1<= rack(0);
      type_cast_863_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_863_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp506x_xop_860,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_53_864,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_883_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_883_inst_req_0;
      type_cast_883_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_883_inst_req_1;
      type_cast_883_inst_ack_1<= rack(0);
      type_cast_883_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_883_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext500_905,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_883_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_88_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_88_inst_req_0;
      type_cast_88_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_88_inst_req_1;
      type_cast_88_inst_ack_1<= rack(0);
      type_cast_88_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_88_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_85,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_89,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_927_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_927_inst_req_0;
      type_cast_927_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_927_inst_req_1;
      type_cast_927_inst_ack_1<= rack(0);
      type_cast_927_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_927_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_926_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv276_928,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1171_index_1_rename
    process(R_indvar_1170_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1170_resized;
      ov(13 downto 0) := iv;
      R_indvar_1170_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1171_index_1_resize
    process(indvar_1159) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1159;
      ov := iv(13 downto 0);
      R_indvar_1170_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1171_root_address_inst
    process(array_obj_ref_1171_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1171_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1171_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_453_index_1_rename
    process(R_indvar529_452_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar529_452_resized;
      ov(13 downto 0) := iv;
      R_indvar529_452_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_453_index_1_resize
    process(indvar529_441) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar529_441;
      ov := iv(13 downto 0);
      R_indvar529_452_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_453_root_address_inst
    process(array_obj_ref_453_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_453_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_453_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_660_index_1_rename
    process(R_indvar513_659_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar513_659_resized;
      ov(10 downto 0) := iv;
      R_indvar513_659_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_660_index_1_resize
    process(indvar513_648) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar513_648;
      ov := iv(10 downto 0);
      R_indvar513_659_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_660_root_address_inst
    process(array_obj_ref_660_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_660_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_660_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_892_index_1_rename
    process(R_indvar499_891_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar499_891_resized;
      ov(13 downto 0) := iv;
      R_indvar499_891_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_892_index_1_resize
    process(indvar499_880) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar499_880;
      ov := iv(13 downto 0);
      R_indvar499_891_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_892_root_address_inst
    process(array_obj_ref_892_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_892_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_892_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1176_addr_0
    process(ptr_deref_1176_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1176_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1176_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1176_base_resize
    process(arrayidx407_1173) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx407_1173;
      ov := iv(13 downto 0);
      ptr_deref_1176_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1176_gather_scatter
    process(ptr_deref_1176_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1176_data_0;
      ov(63 downto 0) := iv;
      tmp408_1177 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1176_root_address_inst
    process(ptr_deref_1176_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1176_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1176_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_590_addr_0
    process(ptr_deref_590_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_590_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_590_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_590_base_resize
    process(arrayidx_455) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_455;
      ov := iv(13 downto 0);
      ptr_deref_590_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_590_gather_scatter
    process(add186_588) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add186_588;
      ov(63 downto 0) := iv;
      ptr_deref_590_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_590_root_address_inst
    process(ptr_deref_590_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_590_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_590_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_797_addr_0
    process(ptr_deref_797_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_797_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_797_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_797_base_resize
    process(arrayidx246_662) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx246_662;
      ov := iv(10 downto 0);
      ptr_deref_797_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_797_gather_scatter
    process(add242_795) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add242_795;
      ov(63 downto 0) := iv;
      ptr_deref_797_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_797_root_address_inst
    process(ptr_deref_797_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_797_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_797_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_896_addr_0
    process(ptr_deref_896_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_896_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_896_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_896_base_resize
    process(arrayidx269_894) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx269_894;
      ov := iv(13 downto 0);
      ptr_deref_896_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_896_gather_scatter
    process(type_cast_898_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_898_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_896_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_896_root_address_inst
    process(ptr_deref_896_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_896_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_896_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1115_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264479_835;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1115_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1115_branch_req_0,
          ack0 => if_stmt_1115_branch_ack_0,
          ack1 => if_stmt_1115_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1287_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1286;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1287_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1287_branch_req_0,
          ack0 => if_stmt_1287_branch_ack_0,
          ack1 => if_stmt_1287_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_388_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp487_387;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_388_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_388_branch_req_0,
          ack0 => if_stmt_388_branch_ack_0,
          ack1 => if_stmt_388_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_403_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp194483_402;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_403_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_403_branch_req_0,
          ack0 => if_stmt_403_branch_ack_0,
          ack1 => if_stmt_403_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_604_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_603;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_604_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_604_branch_req_0,
          ack0 => if_stmt_604_branch_ack_0,
          ack1 => if_stmt_604_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_811_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_810;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_811_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_811_branch_req_0,
          ack0 => if_stmt_811_branch_ack_0,
          ack1 => if_stmt_811_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_836_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp264479_835;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_836_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_836_branch_req_0,
          ack0 => if_stmt_836_branch_ack_0,
          ack1 => if_stmt_836_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_911_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_910;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_911_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_911_branch_req_0,
          ack0 => if_stmt_911_branch_ack_0,
          ack1 => if_stmt_911_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1138_inst
    process(tmp494_1127) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp494_1127, type_cast_1137_wire_constant, tmp_var);
      tmp494x_xop_1139 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_239_inst
    process(add74_235, shr_223) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add74_235, shr_223, tmp_var);
      add79_240 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_420_inst
    process(shr_223) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr_223, type_cast_419_wire_constant, tmp_var);
      tmp536x_xop_421 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_627_inst
    process(tmp522_616) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp522_616, type_cast_626_wire_constant, tmp_var);
      tmp522x_xop_628 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_859_inst
    process(tmp506_848) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp506_848, type_cast_858_wire_constant, tmp_var);
      tmp506x_xop_860 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1148_inst
    process(iNsTr_172_1143) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_172_1143, type_cast_1147_wire_constant, tmp_var);
      xx_xop_1149 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1280_inst
    process(indvar_1159) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1159, type_cast_1279_wire_constant, tmp_var);
      indvarx_xnext_1281 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_430_inst
    process(iNsTr_26_425) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_26_425, type_cast_429_wire_constant, tmp_var);
      xx_xop545_431 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_597_inst
    process(indvar529_441) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar529_441, type_cast_596_wire_constant, tmp_var);
      indvarx_xnext530_598 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_637_inst
    process(iNsTr_39_632) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_39_632, type_cast_636_wire_constant, tmp_var);
      xx_xop544_638 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_804_inst
    process(indvar513_648) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar513_648, type_cast_803_wire_constant, tmp_var);
      indvarx_xnext514_805 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_869_inst
    process(iNsTr_53_864) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_53_864, type_cast_868_wire_constant, tmp_var);
      xx_xop543_870 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_904_inst
    process(indvar499_880) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar499_880, type_cast_903_wire_constant, tmp_var);
      indvarx_xnext500_905 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_234_inst
    process(iNsTr_14_229) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_14_229, type_cast_233_wire_constant, tmp_var);
      add74_235 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1285_inst
    process(indvarx_xnext_1281, tmp498_1156) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1281, tmp498_1156, tmp_var);
      exitcond1_1286 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_602_inst
    process(indvarx_xnext530_598, tmp541_438) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext530_598, tmp541_438, tmp_var);
      exitcond3_603 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_809_inst
    process(indvarx_xnext514_805, tmp527_645) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext514_805, tmp527_645, tmp_var);
      exitcond2_810 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_909_inst
    process(indvarx_xnext500_905, tmp511_877) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext500_905, tmp511_877, tmp_var);
      exitcond_910 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1126_inst
    process(mul259_829) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_829, type_cast_1125_wire_constant, tmp_var);
      tmp494_1127 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_222_inst
    process(mul66_217) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_217, type_cast_221_wire_constant, tmp_var);
      shr_223 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_228_inst
    process(mul66_217) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul66_217, type_cast_227_wire_constant, tmp_var);
      iNsTr_14_229 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_615_inst
    process(mul91_255) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul91_255, type_cast_614_wire_constant, tmp_var);
      tmp522_616 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_847_inst
    process(mul259_829) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul259_829, type_cast_846_wire_constant, tmp_var);
      tmp506_848 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1186_inst
    process(tmp408_1177) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp408_1177, type_cast_1185_wire_constant, tmp_var);
      shr414_1187 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1196_inst
    process(tmp408_1177) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp408_1177, type_cast_1195_wire_constant, tmp_var);
      shr420_1197 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1206_inst
    process(tmp408_1177) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp408_1177, type_cast_1205_wire_constant, tmp_var);
      shr426_1207 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1216_inst
    process(tmp408_1177) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp408_1177, type_cast_1215_wire_constant, tmp_var);
      shr432_1217 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1226_inst
    process(tmp408_1177) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp408_1177, type_cast_1225_wire_constant, tmp_var);
      shr438_1227 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1236_inst
    process(tmp408_1177) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp408_1177, type_cast_1235_wire_constant, tmp_var);
      shr444_1237 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1246_inst
    process(tmp408_1177) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp408_1177, type_cast_1245_wire_constant, tmp_var);
      shr450_1247 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_211_inst
    process(add12_82, add_57) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add12_82, add_57, tmp_var);
      mul_212 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_216_inst
    process(mul_212, add21_107) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_212, add21_107, tmp_var);
      mul66_217 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_244_inst
    process(add39_157, add30_132) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add39_157, add30_132, tmp_var);
      mul85_245 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_249_inst
    process(mul85_245, add48_182) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul85_245, add48_182, tmp_var);
      mul88_250 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_254_inst
    process(mul88_250, add57_207) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul88_250, add57_207, tmp_var);
      mul91_255 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_823_inst
    process(add126_355, add117_330) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add126_355, add117_330, tmp_var);
      mul256_824 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_828_inst
    process(mul256_824, add135_380) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul256_824, add135_380, tmp_var);
      mul259_829 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_106_inst
    process(shl18_95, conv20_102) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_95, conv20_102, tmp_var);
      add21_107 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_131_inst
    process(shl27_120, conv29_127) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_120, conv29_127, tmp_var);
      add30_132 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_156_inst
    process(shl36_145, conv38_152) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_145, conv38_152, tmp_var);
      add39_157 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_181_inst
    process(shl45_170, conv47_177) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_170, conv47_177, tmp_var);
      add48_182 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_206_inst
    process(shl54_195, conv56_202) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_195, conv56_202, tmp_var);
      add57_207 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_279_inst
    process(shl96_268, conv98_275) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl96_268, conv98_275, tmp_var);
      add99_280 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_304_inst
    process(shl105_293, conv107_300) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl105_293, conv107_300, tmp_var);
      add108_305 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_329_inst
    process(shl114_318, conv116_325) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_318, conv116_325, tmp_var);
      add117_330 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_354_inst
    process(shl123_343, conv125_350) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl123_343, conv125_350, tmp_var);
      add126_355 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_379_inst
    process(shl132_368, conv134_375) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_368, conv134_375, tmp_var);
      add135_380 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_56_inst
    process(shl_45, conv3_52) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_45, conv3_52, tmp_var);
      add_57 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_81_inst
    process(shl9_70, conv11_77) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_70, conv11_77, tmp_var);
      add12_82 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_479_inst
    process(shl146_468, conv149_475) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl146_468, conv149_475, tmp_var);
      add150_480 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_497_inst
    process(shl152_486, conv155_493) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl152_486, conv155_493, tmp_var);
      add156_498 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_515_inst
    process(shl158_504, conv161_511) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl158_504, conv161_511, tmp_var);
      add162_516 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_533_inst
    process(shl164_522, conv167_529) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl164_522, conv167_529, tmp_var);
      add168_534 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_551_inst
    process(shl170_540, conv173_547) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl170_540, conv173_547, tmp_var);
      add174_552 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_569_inst
    process(shl176_558, conv179_565) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl176_558, conv179_565, tmp_var);
      add180_570 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_587_inst
    process(shl182_576, conv185_583) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl182_576, conv185_583, tmp_var);
      add186_588 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_686_inst
    process(shl202_675, conv205_682) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl202_675, conv205_682, tmp_var);
      add206_687 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_704_inst
    process(shl208_693, conv211_700) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl208_693, conv211_700, tmp_var);
      add212_705 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_722_inst
    process(shl214_711, conv217_718) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl214_711, conv217_718, tmp_var);
      add218_723 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_740_inst
    process(shl220_729, conv223_736) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl220_729, conv223_736, tmp_var);
      add224_741 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_758_inst
    process(shl226_747, conv229_754) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl226_747, conv229_754, tmp_var);
      add230_759 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_776_inst
    process(shl232_765, conv235_772) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl232_765, conv235_772, tmp_var);
      add236_777 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_794_inst
    process(shl238_783, conv241_790) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl238_783, conv241_790, tmp_var);
      add242_795 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_119_inst
    process(conv26_114) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_114, type_cast_118_wire_constant, tmp_var);
      shl27_120 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_144_inst
    process(conv35_139) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_139, type_cast_143_wire_constant, tmp_var);
      shl36_145 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_169_inst
    process(conv44_164) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_164, type_cast_168_wire_constant, tmp_var);
      shl45_170 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_194_inst
    process(conv53_189) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_189, type_cast_193_wire_constant, tmp_var);
      shl54_195 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_267_inst
    process(conv95_262) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv95_262, type_cast_266_wire_constant, tmp_var);
      shl96_268 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_292_inst
    process(conv104_287) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv104_287, type_cast_291_wire_constant, tmp_var);
      shl105_293 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_317_inst
    process(conv113_312) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv113_312, type_cast_316_wire_constant, tmp_var);
      shl114_318 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_342_inst
    process(conv122_337) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv122_337, type_cast_341_wire_constant, tmp_var);
      shl123_343 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_367_inst
    process(conv131_362) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv131_362, type_cast_366_wire_constant, tmp_var);
      shl132_368 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_44_inst
    process(conv1_39) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_39, type_cast_43_wire_constant, tmp_var);
      shl_45 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_69_inst
    process(conv8_64) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_64, type_cast_68_wire_constant, tmp_var);
      shl9_70 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_94_inst
    process(conv17_89) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_89, type_cast_93_wire_constant, tmp_var);
      shl18_95 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_467_inst
    process(conv144_462) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv144_462, type_cast_466_wire_constant, tmp_var);
      shl146_468 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_485_inst
    process(add150_480) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add150_480, type_cast_484_wire_constant, tmp_var);
      shl152_486 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_503_inst
    process(add156_498) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add156_498, type_cast_502_wire_constant, tmp_var);
      shl158_504 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_521_inst
    process(add162_516) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add162_516, type_cast_520_wire_constant, tmp_var);
      shl164_522 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_539_inst
    process(add168_534) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add168_534, type_cast_538_wire_constant, tmp_var);
      shl170_540 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_557_inst
    process(add174_552) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add174_552, type_cast_556_wire_constant, tmp_var);
      shl176_558 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_575_inst
    process(add180_570) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add180_570, type_cast_574_wire_constant, tmp_var);
      shl182_576 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_674_inst
    process(conv200_669) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv200_669, type_cast_673_wire_constant, tmp_var);
      shl202_675 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_692_inst
    process(add206_687) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add206_687, type_cast_691_wire_constant, tmp_var);
      shl208_693 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_710_inst
    process(add212_705) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add212_705, type_cast_709_wire_constant, tmp_var);
      shl214_711 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_728_inst
    process(add218_723) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add218_723, type_cast_727_wire_constant, tmp_var);
      shl220_729 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_746_inst
    process(add224_741) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add224_741, type_cast_745_wire_constant, tmp_var);
      shl226_747 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_764_inst
    process(add230_759) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add230_759, type_cast_763_wire_constant, tmp_var);
      shl232_765 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_782_inst
    process(add236_777) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add236_777, type_cast_781_wire_constant, tmp_var);
      shl238_783 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1109_inst
    process(conv391_1105, conv276_928) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv391_1105, conv276_928, tmp_var);
      sub_1110 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1132_inst
    process(tmp494_1127) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp494_1127, type_cast_1131_wire_constant, tmp_var);
      tmp495_1133 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_385_inst
    process(mul66_217) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul66_217, type_cast_384_wire_constant, tmp_var);
      cmp487_387 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_401_inst
    process(mul91_255) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul91_255, type_cast_400_wire_constant, tmp_var);
      cmp194483_402 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_414_inst
    process(shr_223) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_223, type_cast_413_wire_constant, tmp_var);
      tmp537_415 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_621_inst
    process(tmp522_616) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp522_616, type_cast_620_wire_constant, tmp_var);
      tmp523_622 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_834_inst
    process(mul259_829) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul259_829, type_cast_833_wire_constant, tmp_var);
      cmp264479_835 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_853_inst
    process(tmp506_848) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp506_848, type_cast_852_wire_constant, tmp_var);
      tmp507_854 <= tmp_var; --
    end process;
    -- shared split operator group (97) : array_obj_ref_1171_index_offset 
    ApIntAdd_group_97: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1170_scaled;
      array_obj_ref_1171_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1171_index_offset_req_0;
      array_obj_ref_1171_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1171_index_offset_req_1;
      array_obj_ref_1171_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_97_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_97_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_97",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 97
    -- shared split operator group (98) : array_obj_ref_453_index_offset 
    ApIntAdd_group_98: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar529_452_scaled;
      array_obj_ref_453_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_453_index_offset_req_0;
      array_obj_ref_453_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_453_index_offset_req_1;
      array_obj_ref_453_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_98_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_98_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_98",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 98
    -- shared split operator group (99) : array_obj_ref_660_index_offset 
    ApIntAdd_group_99: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar513_659_scaled;
      array_obj_ref_660_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_660_index_offset_req_0;
      array_obj_ref_660_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_660_index_offset_req_1;
      array_obj_ref_660_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_99_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_99_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_99",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100010",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 99
    -- shared split operator group (100) : array_obj_ref_892_index_offset 
    ApIntAdd_group_100: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar499_891_scaled;
      array_obj_ref_892_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_892_index_offset_req_0;
      array_obj_ref_892_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_892_index_offset_req_1;
      array_obj_ref_892_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_100_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_100_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_100",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 100
    -- unary operator type_cast_1103_inst
    process(call390_1100) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call390_1100, tmp_var);
      type_cast_1103_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_926_inst
    process(call275_922) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call275_922, tmp_var);
      type_cast_926_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1176_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1176_load_0_req_0;
      ptr_deref_1176_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1176_load_0_req_1;
      ptr_deref_1176_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1176_word_address_0;
      ptr_deref_1176_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_590_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_590_store_0_req_0;
      ptr_deref_590_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_590_store_0_req_1;
      ptr_deref_590_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_590_word_address_0;
      data_in <= ptr_deref_590_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_797_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_797_store_0_req_0;
      ptr_deref_797_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_797_store_0_req_1;
      ptr_deref_797_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_797_word_address_0;
      data_in <= ptr_deref_797_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(10 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_896_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_896_store_0_req_0;
      ptr_deref_896_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_896_store_0_req_1;
      ptr_deref_896_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_896_word_address_0;
      data_in <= ptr_deref_896_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared inport operator group (0) : RPIPE_Block0_done_1087_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1087_inst_req_0;
      RPIPE_Block0_done_1087_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1087_inst_req_1;
      RPIPE_Block0_done_1087_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call378_1088 <= data_out(31 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1090_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1090_inst_req_0;
      RPIPE_Block1_done_1090_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1090_inst_req_1;
      RPIPE_Block1_done_1090_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call381_1091 <= data_out(31 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1093_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1093_inst_req_0;
      RPIPE_Block2_done_1093_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1093_inst_req_1;
      RPIPE_Block2_done_1093_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call384_1094 <= data_out(31 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1096_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1096_inst_req_0;
      RPIPE_Block3_done_1096_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1096_inst_req_1;
      RPIPE_Block3_done_1096_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call387_1097 <= data_out(31 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_ConvTranspose_input_pipe_488_inst RPIPE_ConvTranspose_input_pipe_282_inst RPIPE_ConvTranspose_input_pipe_320_inst RPIPE_ConvTranspose_input_pipe_370_inst RPIPE_ConvTranspose_input_pipe_270_inst RPIPE_ConvTranspose_input_pipe_506_inst RPIPE_ConvTranspose_input_pipe_172_inst RPIPE_ConvTranspose_input_pipe_295_inst RPIPE_ConvTranspose_input_pipe_524_inst RPIPE_ConvTranspose_input_pipe_470_inst RPIPE_ConvTranspose_input_pipe_332_inst RPIPE_ConvTranspose_input_pipe_307_inst RPIPE_ConvTranspose_input_pipe_560_inst RPIPE_ConvTranspose_input_pipe_257_inst RPIPE_ConvTranspose_input_pipe_457_inst RPIPE_ConvTranspose_input_pipe_34_inst RPIPE_ConvTranspose_input_pipe_47_inst RPIPE_ConvTranspose_input_pipe_197_inst RPIPE_ConvTranspose_input_pipe_59_inst RPIPE_ConvTranspose_input_pipe_159_inst RPIPE_ConvTranspose_input_pipe_72_inst RPIPE_ConvTranspose_input_pipe_84_inst RPIPE_ConvTranspose_input_pipe_184_inst RPIPE_ConvTranspose_input_pipe_345_inst RPIPE_ConvTranspose_input_pipe_357_inst RPIPE_ConvTranspose_input_pipe_542_inst RPIPE_ConvTranspose_input_pipe_785_inst RPIPE_ConvTranspose_input_pipe_767_inst RPIPE_ConvTranspose_input_pipe_749_inst RPIPE_ConvTranspose_input_pipe_147_inst RPIPE_ConvTranspose_input_pipe_731_inst RPIPE_ConvTranspose_input_pipe_713_inst RPIPE_ConvTranspose_input_pipe_695_inst RPIPE_ConvTranspose_input_pipe_134_inst RPIPE_ConvTranspose_input_pipe_677_inst RPIPE_ConvTranspose_input_pipe_664_inst RPIPE_ConvTranspose_input_pipe_122_inst RPIPE_ConvTranspose_input_pipe_109_inst RPIPE_ConvTranspose_input_pipe_97_inst RPIPE_ConvTranspose_input_pipe_578_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(319 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 39 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 39 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 39 downto 0);
      signal guard_vector : std_logic_vector( 39 downto 0);
      constant outBUFs : IntegerArray(39 downto 0) := (39 => 1, 38 => 1, 37 => 1, 36 => 1, 35 => 1, 34 => 1, 33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(39 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false, 35 => false, 36 => false, 37 => false, 38 => false, 39 => false);
      constant guardBuffering: IntegerArray(39 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2, 35 => 2, 36 => 2, 37 => 2, 38 => 2, 39 => 2);
      -- 
    begin -- 
      reqL_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_488_inst_req_0;
      reqL_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_282_inst_req_0;
      reqL_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_320_inst_req_0;
      reqL_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_370_inst_req_0;
      reqL_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_270_inst_req_0;
      reqL_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_506_inst_req_0;
      reqL_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_172_inst_req_0;
      reqL_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_295_inst_req_0;
      reqL_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_524_inst_req_0;
      reqL_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_470_inst_req_0;
      reqL_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_332_inst_req_0;
      reqL_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_307_inst_req_0;
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_560_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_257_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_457_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_47_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_197_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_59_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_159_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_72_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_84_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_184_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_345_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_357_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_542_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_785_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_767_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_749_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_147_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_731_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_713_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_695_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_134_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_677_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_664_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_122_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_109_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_97_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_578_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_488_inst_ack_0 <= ackL_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_282_inst_ack_0 <= ackL_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_320_inst_ack_0 <= ackL_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_370_inst_ack_0 <= ackL_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_270_inst_ack_0 <= ackL_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_506_inst_ack_0 <= ackL_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_172_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_295_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_524_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_470_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_332_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_307_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_560_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_257_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_457_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_47_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_197_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_59_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_159_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_72_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_84_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_184_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_345_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_357_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_542_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_785_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_767_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_749_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_147_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_731_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_713_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_695_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_134_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_677_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_664_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_122_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_109_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_97_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_578_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(39) <= RPIPE_ConvTranspose_input_pipe_488_inst_req_1;
      reqR_unguarded(38) <= RPIPE_ConvTranspose_input_pipe_282_inst_req_1;
      reqR_unguarded(37) <= RPIPE_ConvTranspose_input_pipe_320_inst_req_1;
      reqR_unguarded(36) <= RPIPE_ConvTranspose_input_pipe_370_inst_req_1;
      reqR_unguarded(35) <= RPIPE_ConvTranspose_input_pipe_270_inst_req_1;
      reqR_unguarded(34) <= RPIPE_ConvTranspose_input_pipe_506_inst_req_1;
      reqR_unguarded(33) <= RPIPE_ConvTranspose_input_pipe_172_inst_req_1;
      reqR_unguarded(32) <= RPIPE_ConvTranspose_input_pipe_295_inst_req_1;
      reqR_unguarded(31) <= RPIPE_ConvTranspose_input_pipe_524_inst_req_1;
      reqR_unguarded(30) <= RPIPE_ConvTranspose_input_pipe_470_inst_req_1;
      reqR_unguarded(29) <= RPIPE_ConvTranspose_input_pipe_332_inst_req_1;
      reqR_unguarded(28) <= RPIPE_ConvTranspose_input_pipe_307_inst_req_1;
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_560_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_257_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_457_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_47_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_197_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_59_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_159_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_72_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_84_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_184_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_345_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_357_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_542_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_785_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_767_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_749_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_147_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_731_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_713_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_695_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_134_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_677_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_664_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_122_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_109_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_97_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_578_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_488_inst_ack_1 <= ackR_unguarded(39);
      RPIPE_ConvTranspose_input_pipe_282_inst_ack_1 <= ackR_unguarded(38);
      RPIPE_ConvTranspose_input_pipe_320_inst_ack_1 <= ackR_unguarded(37);
      RPIPE_ConvTranspose_input_pipe_370_inst_ack_1 <= ackR_unguarded(36);
      RPIPE_ConvTranspose_input_pipe_270_inst_ack_1 <= ackR_unguarded(35);
      RPIPE_ConvTranspose_input_pipe_506_inst_ack_1 <= ackR_unguarded(34);
      RPIPE_ConvTranspose_input_pipe_172_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_ConvTranspose_input_pipe_295_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_ConvTranspose_input_pipe_524_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_ConvTranspose_input_pipe_470_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_ConvTranspose_input_pipe_332_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_ConvTranspose_input_pipe_307_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_ConvTranspose_input_pipe_560_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_257_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_457_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_47_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_197_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_59_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_159_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_72_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_84_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_184_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_345_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_357_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_542_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_785_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_767_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_749_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_147_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_731_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_713_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_695_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_134_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_677_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_664_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_122_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_109_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_97_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_578_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      guard_vector(35)  <=  '1';
      guard_vector(36)  <=  '1';
      guard_vector(37)  <=  '1';
      guard_vector(38)  <=  '1';
      guard_vector(39)  <=  '1';
      call153_489 <= data_out(319 downto 312);
      call101_283 <= data_out(311 downto 304);
      call115_321 <= data_out(303 downto 296);
      call133_371 <= data_out(295 downto 288);
      call97_271 <= data_out(287 downto 280);
      call159_507 <= data_out(279 downto 272);
      call46_173 <= data_out(271 downto 264);
      call106_296 <= data_out(263 downto 256);
      call165_525 <= data_out(255 downto 248);
      call147_471 <= data_out(247 downto 240);
      call119_333 <= data_out(239 downto 232);
      call110_308 <= data_out(231 downto 224);
      call177_561 <= data_out(223 downto 216);
      call92_258 <= data_out(215 downto 208);
      call143_458 <= data_out(207 downto 200);
      call_35 <= data_out(199 downto 192);
      call2_48 <= data_out(191 downto 184);
      call55_198 <= data_out(183 downto 176);
      call5_60 <= data_out(175 downto 168);
      call41_160 <= data_out(167 downto 160);
      call10_73 <= data_out(159 downto 152);
      call14_85 <= data_out(151 downto 144);
      call50_185 <= data_out(143 downto 136);
      call124_346 <= data_out(135 downto 128);
      call128_358 <= data_out(127 downto 120);
      call171_543 <= data_out(119 downto 112);
      call239_786 <= data_out(111 downto 104);
      call233_768 <= data_out(103 downto 96);
      call227_750 <= data_out(95 downto 88);
      call37_148 <= data_out(87 downto 80);
      call221_732 <= data_out(79 downto 72);
      call215_714 <= data_out(71 downto 64);
      call209_696 <= data_out(63 downto 56);
      call32_135 <= data_out(55 downto 48);
      call203_678 <= data_out(47 downto 40);
      call199_665 <= data_out(39 downto 32);
      call28_123 <= data_out(31 downto 24);
      call23_110 <= data_out(23 downto 16);
      call19_98 <= data_out(15 downto 8);
      call183_579 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_4_gI", nreqs => 40, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_4: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_4", data_width => 8,  num_reqs => 40,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared outport operator group (0) : WPIPE_Block0_start_929_inst WPIPE_Block0_start_932_inst WPIPE_Block0_start_935_inst WPIPE_Block0_start_938_inst WPIPE_Block0_start_941_inst WPIPE_Block0_start_944_inst WPIPE_Block0_start_947_inst WPIPE_Block0_start_950_inst WPIPE_Block0_start_953_inst WPIPE_Block0_start_956_inst WPIPE_Block0_start_960_inst WPIPE_Block0_start_963_inst WPIPE_Block0_start_966_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(415 downto 0);
      signal sample_req, sample_ack : BooleanArray( 12 downto 0);
      signal update_req, update_ack : BooleanArray( 12 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 12 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 12 downto 0);
      signal guard_vector : std_logic_vector( 12 downto 0);
      constant inBUFs : IntegerArray(12 downto 0) := (12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(12 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false);
      constant guardBuffering: IntegerArray(12 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2);
      -- 
    begin -- 
      sample_req_unguarded(12) <= WPIPE_Block0_start_929_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block0_start_932_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block0_start_935_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block0_start_938_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block0_start_941_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block0_start_944_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block0_start_947_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_start_950_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_start_953_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_start_956_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_start_960_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_start_963_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_start_966_inst_req_0;
      WPIPE_Block0_start_929_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block0_start_932_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block0_start_935_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block0_start_938_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block0_start_941_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block0_start_944_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block0_start_947_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_start_950_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_start_953_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_start_956_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_start_960_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_start_963_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_start_966_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(12) <= WPIPE_Block0_start_929_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block0_start_932_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block0_start_935_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block0_start_938_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block0_start_941_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block0_start_944_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block0_start_947_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_start_950_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_start_953_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_start_956_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_start_960_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_start_963_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_start_966_inst_req_1;
      WPIPE_Block0_start_929_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block0_start_932_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block0_start_935_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block0_start_938_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block0_start_941_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block0_start_944_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block0_start_947_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_start_950_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_start_953_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_start_956_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_start_960_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_start_963_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_start_966_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      data_in <= add_57 & add12_82 & add21_107 & add30_132 & add39_157 & add48_182 & add57_207 & add99_280 & add108_305 & type_cast_958_wire_constant & add117_330 & add126_355 & add135_380;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 13, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 32, num_reqs => 13, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_969_inst WPIPE_Block1_start_972_inst WPIPE_Block1_start_975_inst WPIPE_Block1_start_978_inst WPIPE_Block1_start_981_inst WPIPE_Block1_start_984_inst WPIPE_Block1_start_987_inst WPIPE_Block1_start_990_inst WPIPE_Block1_start_993_inst WPIPE_Block1_start_996_inst WPIPE_Block1_start_999_inst WPIPE_Block1_start_1002_inst WPIPE_Block1_start_1005_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(415 downto 0);
      signal sample_req, sample_ack : BooleanArray( 12 downto 0);
      signal update_req, update_ack : BooleanArray( 12 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 12 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 12 downto 0);
      signal guard_vector : std_logic_vector( 12 downto 0);
      constant inBUFs : IntegerArray(12 downto 0) := (12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(12 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false);
      constant guardBuffering: IntegerArray(12 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2);
      -- 
    begin -- 
      sample_req_unguarded(12) <= WPIPE_Block1_start_969_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block1_start_972_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block1_start_975_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block1_start_978_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block1_start_981_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block1_start_984_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block1_start_987_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block1_start_990_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block1_start_993_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block1_start_996_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block1_start_999_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block1_start_1002_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block1_start_1005_inst_req_0;
      WPIPE_Block1_start_969_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block1_start_972_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block1_start_975_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block1_start_978_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block1_start_981_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block1_start_984_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block1_start_987_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block1_start_990_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block1_start_993_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block1_start_996_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block1_start_999_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block1_start_1002_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block1_start_1005_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(12) <= WPIPE_Block1_start_969_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block1_start_972_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block1_start_975_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block1_start_978_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block1_start_981_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block1_start_984_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block1_start_987_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block1_start_990_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block1_start_993_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block1_start_996_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block1_start_999_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block1_start_1002_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block1_start_1005_inst_req_1;
      WPIPE_Block1_start_969_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block1_start_972_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block1_start_975_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block1_start_978_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block1_start_981_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block1_start_984_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block1_start_987_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block1_start_990_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block1_start_993_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block1_start_996_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block1_start_999_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block1_start_1002_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block1_start_1005_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      data_in <= add_57 & add12_82 & add21_107 & add30_132 & add39_157 & add48_182 & add57_207 & add99_280 & add108_305 & shr_223 & add117_330 & add126_355 & add135_380;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 13, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 32, num_reqs => 13, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1008_inst WPIPE_Block2_start_1011_inst WPIPE_Block2_start_1014_inst WPIPE_Block2_start_1017_inst WPIPE_Block2_start_1020_inst WPIPE_Block2_start_1023_inst WPIPE_Block2_start_1026_inst WPIPE_Block2_start_1029_inst WPIPE_Block2_start_1032_inst WPIPE_Block2_start_1035_inst WPIPE_Block2_start_1038_inst WPIPE_Block2_start_1041_inst WPIPE_Block2_start_1044_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(415 downto 0);
      signal sample_req, sample_ack : BooleanArray( 12 downto 0);
      signal update_req, update_ack : BooleanArray( 12 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 12 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 12 downto 0);
      signal guard_vector : std_logic_vector( 12 downto 0);
      constant inBUFs : IntegerArray(12 downto 0) := (12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(12 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false);
      constant guardBuffering: IntegerArray(12 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2);
      -- 
    begin -- 
      sample_req_unguarded(12) <= WPIPE_Block2_start_1008_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block2_start_1011_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block2_start_1014_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block2_start_1017_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block2_start_1020_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block2_start_1023_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block2_start_1026_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block2_start_1029_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block2_start_1032_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block2_start_1035_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block2_start_1038_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block2_start_1041_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block2_start_1044_inst_req_0;
      WPIPE_Block2_start_1008_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block2_start_1011_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block2_start_1014_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block2_start_1017_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block2_start_1020_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block2_start_1023_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block2_start_1026_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block2_start_1029_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block2_start_1032_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block2_start_1035_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block2_start_1038_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block2_start_1041_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block2_start_1044_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(12) <= WPIPE_Block2_start_1008_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block2_start_1011_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block2_start_1014_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block2_start_1017_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block2_start_1020_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block2_start_1023_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block2_start_1026_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block2_start_1029_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block2_start_1032_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block2_start_1035_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block2_start_1038_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block2_start_1041_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block2_start_1044_inst_req_1;
      WPIPE_Block2_start_1008_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block2_start_1011_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block2_start_1014_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block2_start_1017_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block2_start_1020_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block2_start_1023_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block2_start_1026_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block2_start_1029_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block2_start_1032_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block2_start_1035_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block2_start_1038_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block2_start_1041_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block2_start_1044_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      data_in <= add_57 & add12_82 & add21_107 & add30_132 & add39_157 & add48_182 & add57_207 & add99_280 & add108_305 & add74_235 & add117_330 & add126_355 & add135_380;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 13, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 32, num_reqs => 13, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1047_inst WPIPE_Block3_start_1050_inst WPIPE_Block3_start_1053_inst WPIPE_Block3_start_1056_inst WPIPE_Block3_start_1059_inst WPIPE_Block3_start_1062_inst WPIPE_Block3_start_1065_inst WPIPE_Block3_start_1068_inst WPIPE_Block3_start_1071_inst WPIPE_Block3_start_1074_inst WPIPE_Block3_start_1077_inst WPIPE_Block3_start_1080_inst WPIPE_Block3_start_1083_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(415 downto 0);
      signal sample_req, sample_ack : BooleanArray( 12 downto 0);
      signal update_req, update_ack : BooleanArray( 12 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 12 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 12 downto 0);
      signal guard_vector : std_logic_vector( 12 downto 0);
      constant inBUFs : IntegerArray(12 downto 0) := (12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(12 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false);
      constant guardBuffering: IntegerArray(12 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2);
      -- 
    begin -- 
      sample_req_unguarded(12) <= WPIPE_Block3_start_1047_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Block3_start_1050_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Block3_start_1053_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Block3_start_1056_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Block3_start_1059_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Block3_start_1062_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Block3_start_1065_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block3_start_1068_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block3_start_1071_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block3_start_1074_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block3_start_1077_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block3_start_1080_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block3_start_1083_inst_req_0;
      WPIPE_Block3_start_1047_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Block3_start_1050_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Block3_start_1053_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Block3_start_1056_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Block3_start_1059_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Block3_start_1062_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Block3_start_1065_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block3_start_1068_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block3_start_1071_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block3_start_1074_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block3_start_1077_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block3_start_1080_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block3_start_1083_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(12) <= WPIPE_Block3_start_1047_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Block3_start_1050_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Block3_start_1053_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Block3_start_1056_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Block3_start_1059_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Block3_start_1062_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Block3_start_1065_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block3_start_1068_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block3_start_1071_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block3_start_1074_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block3_start_1077_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block3_start_1080_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block3_start_1083_inst_req_1;
      WPIPE_Block3_start_1047_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Block3_start_1050_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Block3_start_1053_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Block3_start_1056_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Block3_start_1059_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Block3_start_1062_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Block3_start_1065_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block3_start_1068_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block3_start_1071_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block3_start_1074_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block3_start_1077_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block3_start_1080_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block3_start_1083_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      data_in <= add_57 & add12_82 & add21_107 & add30_132 & add39_157 & add48_182 & add57_207 & add99_280 & add108_305 & add79_240 & add117_330 & add126_355 & add135_380;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 13, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 32, num_reqs => 13, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_ConvTranspose_output_pipe_1252_inst WPIPE_ConvTranspose_output_pipe_1255_inst WPIPE_ConvTranspose_output_pipe_1258_inst WPIPE_ConvTranspose_output_pipe_1261_inst WPIPE_ConvTranspose_output_pipe_1264_inst WPIPE_ConvTranspose_output_pipe_1267_inst WPIPE_ConvTranspose_output_pipe_1270_inst WPIPE_ConvTranspose_output_pipe_1273_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1252_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1255_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1258_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1261_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1264_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1267_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1270_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1273_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1252_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1255_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1258_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1261_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1264_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1267_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1270_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1273_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1252_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1255_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1258_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1261_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1264_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1267_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1270_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1273_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1252_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1255_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1258_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1261_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1264_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1267_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1270_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1273_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv453_1251 & conv447_1241 & conv441_1231 & conv435_1221 & conv429_1211 & conv423_1201 & conv417_1191 & conv411_1181;
      ConvTranspose_output_pipe_write_4_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_4_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared outport operator group (5) : WPIPE_elapsed_time_pipe_1111_inst 
    OutportGroup_5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1111_inst_req_0;
      WPIPE_elapsed_time_pipe_1111_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1111_inst_req_1;
      WPIPE_elapsed_time_pipe_1111_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub_1110;
      elapsed_time_pipe_write_5_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_5: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- shared call operator group (0) : call_stmt_922_call call_stmt_1100_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_922_call_req_0;
      reqL_unguarded(0) <= call_stmt_1100_call_req_0;
      call_stmt_922_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1100_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_922_call_req_1;
      reqR_unguarded(0) <= call_stmt_1100_call_req_1;
      call_stmt_922_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1100_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call275_922 <= data_out(127 downto 64);
      call390_1100 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(31 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3268_start: Boolean;
  signal convTransposeA_CP_3268_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block0_start_1318_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1330_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1303_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1303_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1306_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1333_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1309_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1336_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1336_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1312_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1339_inst_ack_0 : boolean;
  signal type_cast_1638_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1312_inst_req_1 : boolean;
  signal type_cast_1465_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1306_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1306_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1312_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1339_inst_ack_1 : boolean;
  signal type_cast_1465_inst_ack_0 : boolean;
  signal phi_stmt_1641_ack_0 : boolean;
  signal type_cast_1465_inst_req_0 : boolean;
  signal type_cast_1451_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1312_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1309_inst_req_1 : boolean;
  signal phi_stmt_1628_ack_0 : boolean;
  signal RPIPE_Block0_start_1333_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1330_inst_ack_1 : boolean;
  signal phi_stmt_1635_ack_0 : boolean;
  signal RPIPE_Block0_start_1303_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1321_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1321_inst_req_1 : boolean;
  signal phi_stmt_1628_req_0 : boolean;
  signal RPIPE_Block0_start_1306_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1336_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1321_inst_req_0 : boolean;
  signal type_cast_1465_inst_ack_1 : boolean;
  signal type_cast_1521_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1336_inst_ack_1 : boolean;
  signal type_cast_1479_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1324_inst_req_0 : boolean;
  signal type_cast_1479_inst_ack_0 : boolean;
  signal type_cast_1451_inst_req_1 : boolean;
  signal type_cast_1479_inst_req_1 : boolean;
  signal type_cast_1479_inst_ack_1 : boolean;
  signal type_cast_1451_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1324_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1315_inst_req_0 : boolean;
  signal phi_stmt_1635_req_0 : boolean;
  signal type_cast_1638_inst_req_0 : boolean;
  signal type_cast_1638_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1315_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1339_inst_req_1 : boolean;
  signal type_cast_1521_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1333_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1315_inst_req_1 : boolean;
  signal type_cast_1521_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1330_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1315_inst_ack_1 : boolean;
  signal type_cast_1638_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1318_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1303_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1309_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1333_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1330_inst_ack_0 : boolean;
  signal type_cast_1521_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1309_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1318_inst_ack_1 : boolean;
  signal RPIPE_Block0_start_1318_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1339_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1321_inst_ack_0 : boolean;
  signal type_cast_1451_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1324_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1327_inst_ack_1 : boolean;
  signal type_cast_1646_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1327_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1327_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1327_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1324_inst_ack_1 : boolean;
  signal type_cast_1646_inst_ack_0 : boolean;
  signal type_cast_1640_inst_req_1 : boolean;
  signal array_obj_ref_1527_index_offset_req_0 : boolean;
  signal array_obj_ref_1527_index_offset_ack_0 : boolean;
  signal array_obj_ref_1527_index_offset_req_1 : boolean;
  signal array_obj_ref_1527_index_offset_ack_1 : boolean;
  signal addr_of_1528_final_reg_req_0 : boolean;
  signal addr_of_1528_final_reg_ack_0 : boolean;
  signal phi_stmt_1641_req_0 : boolean;
  signal addr_of_1528_final_reg_req_1 : boolean;
  signal addr_of_1528_final_reg_ack_1 : boolean;
  signal type_cast_1644_inst_ack_1 : boolean;
  signal ptr_deref_1532_load_0_req_0 : boolean;
  signal ptr_deref_1532_load_0_ack_0 : boolean;
  signal phi_stmt_1641_req_1 : boolean;
  signal ptr_deref_1532_load_0_req_1 : boolean;
  signal ptr_deref_1532_load_0_ack_1 : boolean;
  signal phi_stmt_1628_req_1 : boolean;
  signal type_cast_1542_inst_req_0 : boolean;
  signal type_cast_1542_inst_ack_0 : boolean;
  signal type_cast_1644_inst_req_1 : boolean;
  signal type_cast_1542_inst_req_1 : boolean;
  signal type_cast_1542_inst_ack_1 : boolean;
  signal type_cast_1634_inst_ack_1 : boolean;
  signal type_cast_1634_inst_req_1 : boolean;
  signal array_obj_ref_1548_index_offset_req_0 : boolean;
  signal array_obj_ref_1548_index_offset_ack_0 : boolean;
  signal array_obj_ref_1548_index_offset_req_1 : boolean;
  signal array_obj_ref_1548_index_offset_ack_1 : boolean;
  signal type_cast_1634_inst_ack_0 : boolean;
  signal phi_stmt_1635_req_1 : boolean;
  signal addr_of_1549_final_reg_req_0 : boolean;
  signal addr_of_1549_final_reg_ack_0 : boolean;
  signal type_cast_1644_inst_ack_0 : boolean;
  signal addr_of_1549_final_reg_req_1 : boolean;
  signal addr_of_1549_final_reg_ack_1 : boolean;
  signal type_cast_1634_inst_req_0 : boolean;
  signal type_cast_1644_inst_req_0 : boolean;
  signal type_cast_1646_inst_ack_1 : boolean;
  signal type_cast_1646_inst_req_1 : boolean;
  signal ptr_deref_1552_store_0_req_0 : boolean;
  signal ptr_deref_1552_store_0_ack_0 : boolean;
  signal ptr_deref_1552_store_0_req_1 : boolean;
  signal ptr_deref_1552_store_0_ack_1 : boolean;
  signal type_cast_1640_inst_ack_1 : boolean;
  signal type_cast_1640_inst_ack_0 : boolean;
  signal if_stmt_1566_branch_req_0 : boolean;
  signal type_cast_1640_inst_req_0 : boolean;
  signal if_stmt_1566_branch_ack_1 : boolean;
  signal if_stmt_1566_branch_ack_0 : boolean;
  signal type_cast_1589_inst_req_0 : boolean;
  signal type_cast_1589_inst_ack_0 : boolean;
  signal type_cast_1589_inst_req_1 : boolean;
  signal type_cast_1589_inst_ack_1 : boolean;
  signal type_cast_1598_inst_req_0 : boolean;
  signal type_cast_1598_inst_ack_0 : boolean;
  signal type_cast_1598_inst_req_1 : boolean;
  signal type_cast_1598_inst_ack_1 : boolean;
  signal type_cast_1614_inst_req_0 : boolean;
  signal type_cast_1614_inst_ack_0 : boolean;
  signal type_cast_1614_inst_req_1 : boolean;
  signal type_cast_1614_inst_ack_1 : boolean;
  signal if_stmt_1621_branch_req_0 : boolean;
  signal if_stmt_1621_branch_ack_1 : boolean;
  signal if_stmt_1621_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1657_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1657_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1657_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1657_inst_ack_1 : boolean;
  signal phi_stmt_1408_req_0 : boolean;
  signal phi_stmt_1415_req_0 : boolean;
  signal phi_stmt_1423_req_0 : boolean;
  signal phi_stmt_1430_req_0 : boolean;
  signal type_cast_1414_inst_req_0 : boolean;
  signal type_cast_1414_inst_ack_0 : boolean;
  signal type_cast_1414_inst_req_1 : boolean;
  signal type_cast_1414_inst_ack_1 : boolean;
  signal phi_stmt_1408_req_1 : boolean;
  signal type_cast_1422_inst_req_0 : boolean;
  signal type_cast_1422_inst_ack_0 : boolean;
  signal type_cast_1422_inst_req_1 : boolean;
  signal type_cast_1422_inst_ack_1 : boolean;
  signal phi_stmt_1415_req_1 : boolean;
  signal type_cast_1429_inst_req_0 : boolean;
  signal type_cast_1429_inst_ack_0 : boolean;
  signal type_cast_1429_inst_req_1 : boolean;
  signal type_cast_1429_inst_ack_1 : boolean;
  signal phi_stmt_1423_req_1 : boolean;
  signal type_cast_1436_inst_req_0 : boolean;
  signal type_cast_1436_inst_ack_0 : boolean;
  signal type_cast_1436_inst_req_1 : boolean;
  signal type_cast_1436_inst_ack_1 : boolean;
  signal phi_stmt_1430_req_1 : boolean;
  signal phi_stmt_1408_ack_0 : boolean;
  signal phi_stmt_1415_ack_0 : boolean;
  signal phi_stmt_1423_ack_0 : boolean;
  signal phi_stmt_1430_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3268_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3268_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3268_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3268_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3268: Block -- control-path 
    signal convTransposeA_CP_3268_elements: BooleanArray(111 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3268_elements(0) <= convTransposeA_CP_3268_start;
    convTransposeA_CP_3268_symbol <= convTransposeA_CP_3268_elements(64);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340__entry__
      -- CP-element group 0: 	 branch_block_stmt_1301/$entry
      -- CP-element group 0: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1303_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1303_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/$entry
      -- CP-element group 0: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1303_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1301/branch_block_stmt_1301__entry__
      -- CP-element group 0: 	 $entry
      -- 
    rr_3316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(0), ack => RPIPE_Block0_start_1303_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	111 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	70 
    -- CP-element group 1: 	71 
    -- CP-element group 1: 	73 
    -- CP-element group 1: 	74 
    -- CP-element group 1: 	76 
    -- CP-element group 1: 	77 
    -- CP-element group 1: 	79 
    -- CP-element group 1: 	80 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1301/merge_stmt_1627__exit__
      -- CP-element group 1: 	 branch_block_stmt_1301/assign_stmt_1653__entry__
      -- CP-element group 1: 	 branch_block_stmt_1301/assign_stmt_1653__exit__
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1301/assign_stmt_1653/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/assign_stmt_1653/$exit
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1408/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1414/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1414/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1414/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1414/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1414/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1414/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1415/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_sources/type_cast_1422/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_sources/type_cast_1422/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_sources/type_cast_1422/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_sources/type_cast_1422/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_sources/type_cast_1422/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_sources/type_cast_1422/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1423/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1430/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_sources/type_cast_1436/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_sources/type_cast_1436/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_sources/type_cast_1436/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_sources/type_cast_1436/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_sources/type_cast_1436/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_sources/type_cast_1436/SplitProtocol/Update/cr
      -- 
    rr_3918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(1), ack => type_cast_1414_inst_req_0); -- 
    cr_3923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(1), ack => type_cast_1414_inst_req_1); -- 
    rr_3941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(1), ack => type_cast_1422_inst_req_0); -- 
    cr_3946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(1), ack => type_cast_1422_inst_req_1); -- 
    rr_3964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(1), ack => type_cast_1429_inst_req_0); -- 
    cr_3969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(1), ack => type_cast_1429_inst_req_1); -- 
    rr_3987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(1), ack => type_cast_1436_inst_req_0); -- 
    cr_3992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(1), ack => type_cast_1436_inst_req_1); -- 
    convTransposeA_CP_3268_elements(1) <= convTransposeA_CP_3268_elements(111);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1303_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1303_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1303_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1303_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1303_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1303_Sample/$exit
      -- 
    ra_3317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1303_inst_ack_0, ack => convTransposeA_CP_3268_elements(2)); -- 
    cr_3321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(2), ack => RPIPE_Block0_start_1303_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1303_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1306_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1306_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1303_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1306_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1303_update_completed_
      -- 
    ca_3322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1303_inst_ack_1, ack => convTransposeA_CP_3268_elements(3)); -- 
    rr_3330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(3), ack => RPIPE_Block0_start_1306_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1306_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1306_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1306_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1306_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1306_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1306_sample_completed_
      -- 
    ra_3331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1306_inst_ack_0, ack => convTransposeA_CP_3268_elements(4)); -- 
    cr_3335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(4), ack => RPIPE_Block0_start_1306_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1306_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1306_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1306_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1309_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1309_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1309_Sample/rr
      -- 
    ca_3336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1306_inst_ack_1, ack => convTransposeA_CP_3268_elements(5)); -- 
    rr_3344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(5), ack => RPIPE_Block0_start_1309_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1309_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1309_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1309_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1309_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1309_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1309_Sample/ra
      -- 
    ra_3345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1309_inst_ack_0, ack => convTransposeA_CP_3268_elements(6)); -- 
    cr_3349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(6), ack => RPIPE_Block0_start_1309_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1312_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1309_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1312_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1312_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1309_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1309_update_completed_
      -- 
    ca_3350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1309_inst_ack_1, ack => convTransposeA_CP_3268_elements(7)); -- 
    rr_3358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(7), ack => RPIPE_Block0_start_1312_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1312_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1312_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1312_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1312_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1312_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1312_update_start_
      -- 
    ra_3359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1312_inst_ack_0, ack => convTransposeA_CP_3268_elements(8)); -- 
    cr_3363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(8), ack => RPIPE_Block0_start_1312_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1312_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1315_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1312_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1312_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1315_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1315_Sample/rr
      -- 
    ca_3364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1312_inst_ack_1, ack => convTransposeA_CP_3268_elements(9)); -- 
    rr_3372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(9), ack => RPIPE_Block0_start_1315_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1315_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1315_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1315_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1315_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1315_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1315_Update/cr
      -- 
    ra_3373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1315_inst_ack_0, ack => convTransposeA_CP_3268_elements(10)); -- 
    cr_3377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(10), ack => RPIPE_Block0_start_1315_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1315_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1315_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1315_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1318_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1318_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1318_Sample/rr
      -- 
    ca_3378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1315_inst_ack_1, ack => convTransposeA_CP_3268_elements(11)); -- 
    rr_3386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(11), ack => RPIPE_Block0_start_1318_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1318_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1318_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1318_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1318_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1318_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1318_Sample/$exit
      -- 
    ra_3387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1318_inst_ack_0, ack => convTransposeA_CP_3268_elements(12)); -- 
    cr_3391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(12), ack => RPIPE_Block0_start_1318_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1321_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1321_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1318_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1318_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1318_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1321_sample_start_
      -- 
    ca_3392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1318_inst_ack_1, ack => convTransposeA_CP_3268_elements(13)); -- 
    rr_3400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(13), ack => RPIPE_Block0_start_1321_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1321_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1321_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1321_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1321_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1321_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1321_Sample/ra
      -- 
    ra_3401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1321_inst_ack_0, ack => convTransposeA_CP_3268_elements(14)); -- 
    cr_3405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(14), ack => RPIPE_Block0_start_1321_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1321_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1321_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1324_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1324_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1321_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1324_Sample/rr
      -- 
    ca_3406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1321_inst_ack_1, ack => convTransposeA_CP_3268_elements(15)); -- 
    rr_3414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(15), ack => RPIPE_Block0_start_1324_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1324_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1324_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1324_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1324_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1324_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1324_Update/cr
      -- 
    ra_3415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1324_inst_ack_0, ack => convTransposeA_CP_3268_elements(16)); -- 
    cr_3419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(16), ack => RPIPE_Block0_start_1324_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1324_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1324_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1327_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1327_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1327_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1324_Update/ca
      -- 
    ca_3420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1324_inst_ack_1, ack => convTransposeA_CP_3268_elements(17)); -- 
    rr_3428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(17), ack => RPIPE_Block0_start_1327_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1327_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1327_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1327_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1327_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1327_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1327_Sample/$exit
      -- 
    ra_3429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1327_inst_ack_0, ack => convTransposeA_CP_3268_elements(18)); -- 
    cr_3433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(18), ack => RPIPE_Block0_start_1327_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1330_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1330_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1330_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1327_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1327_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1327_Update/$exit
      -- 
    ca_3434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1327_inst_ack_1, ack => convTransposeA_CP_3268_elements(19)); -- 
    rr_3442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(19), ack => RPIPE_Block0_start_1330_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1330_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1330_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1330_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1330_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1330_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1330_update_start_
      -- 
    ra_3443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1330_inst_ack_0, ack => convTransposeA_CP_3268_elements(20)); -- 
    cr_3447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(20), ack => RPIPE_Block0_start_1330_inst_req_1); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1330_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1333_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1330_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1333_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1333_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1330_update_completed_
      -- 
    ca_3448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1330_inst_ack_1, ack => convTransposeA_CP_3268_elements(21)); -- 
    rr_3456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(21), ack => RPIPE_Block0_start_1333_inst_req_0); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1333_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1333_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1333_Update/cr
      -- CP-element group 22: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1333_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1333_update_start_
      -- CP-element group 22: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1333_Update/$entry
      -- 
    ra_3457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1333_inst_ack_0, ack => convTransposeA_CP_3268_elements(22)); -- 
    cr_3461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(22), ack => RPIPE_Block0_start_1333_inst_req_1); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1336_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1336_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1336_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1333_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1333_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1333_update_completed_
      -- 
    ca_3462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1333_inst_ack_1, ack => convTransposeA_CP_3268_elements(23)); -- 
    rr_3470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(23), ack => RPIPE_Block0_start_1336_inst_req_0); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1336_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1336_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1336_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1336_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1336_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1336_Sample/ra
      -- 
    ra_3471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1336_inst_ack_0, ack => convTransposeA_CP_3268_elements(24)); -- 
    cr_3475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(24), ack => RPIPE_Block0_start_1336_inst_req_1); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1336_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1339_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1336_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1336_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1339_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1339_Sample/rr
      -- 
    ca_3476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1336_inst_ack_1, ack => convTransposeA_CP_3268_elements(25)); -- 
    rr_3484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(25), ack => RPIPE_Block0_start_1339_inst_req_0); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1339_update_start_
      -- CP-element group 26: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1339_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1339_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1339_Update/cr
      -- CP-element group 26: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1339_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1339_Sample/$exit
      -- 
    ra_3485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1339_inst_ack_0, ack => convTransposeA_CP_3268_elements(26)); -- 
    cr_3489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(26), ack => RPIPE_Block0_start_1339_inst_req_1); -- 
    -- CP-element group 27:  fork  transition  place  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	65 
    -- CP-element group 27: 	66 
    -- CP-element group 27: 	67 
    -- CP-element group 27: 	68 
    -- CP-element group 27:  members (19) 
      -- CP-element group 27: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340__exit__
      -- CP-element group 27: 	 branch_block_stmt_1301/assign_stmt_1347_to_assign_stmt_1405__entry__
      -- CP-element group 27: 	 branch_block_stmt_1301/entry_whilex_xbody
      -- CP-element group 27: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1339_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1301/assign_stmt_1347_to_assign_stmt_1405__exit__
      -- CP-element group 27: 	 branch_block_stmt_1301/assign_stmt_1347_to_assign_stmt_1405/$entry
      -- CP-element group 27: 	 branch_block_stmt_1301/assign_stmt_1347_to_assign_stmt_1405/$exit
      -- CP-element group 27: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1339_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/RPIPE_Block0_start_1339_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1301/assign_stmt_1304_to_assign_stmt_1340/$exit
      -- CP-element group 27: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 27: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1408/$entry
      -- CP-element group 27: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/$entry
      -- CP-element group 27: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1415/$entry
      -- CP-element group 27: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_sources/$entry
      -- CP-element group 27: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1423/$entry
      -- CP-element group 27: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/$entry
      -- CP-element group 27: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1430/$entry
      -- CP-element group 27: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_sources/$entry
      -- 
    ca_3490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1339_inst_ack_1, ack => convTransposeA_CP_3268_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	88 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1451_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1451_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1451_sample_completed_
      -- 
    ra_3505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1451_inst_ack_0, ack => convTransposeA_CP_3268_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	88 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	42 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1451_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1451_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1451_update_completed_
      -- 
    ca_3510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1451_inst_ack_1, ack => convTransposeA_CP_3268_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	88 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1465_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1465_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1465_Sample/$exit
      -- 
    ra_3519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1465_inst_ack_0, ack => convTransposeA_CP_3268_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	88 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	42 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1465_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1465_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1465_update_completed_
      -- 
    ca_3524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1465_inst_ack_1, ack => convTransposeA_CP_3268_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	88 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1479_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1479_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1479_Sample/$exit
      -- 
    ra_3533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1479_inst_ack_0, ack => convTransposeA_CP_3268_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	88 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	42 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1479_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1479_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1479_update_completed_
      -- 
    ca_3538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1479_inst_ack_1, ack => convTransposeA_CP_3268_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	88 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1521_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1521_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1521_Sample/ra
      -- 
    ra_3547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1521_inst_ack_0, ack => convTransposeA_CP_3268_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	88 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (16) 
      -- CP-element group 35: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_index_resized_1
      -- CP-element group 35: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1521_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_index_scaled_1
      -- CP-element group 35: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_index_computed_1
      -- CP-element group 35: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1521_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1521_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_index_resize_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_index_resize_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_index_resize_1/index_resize_req
      -- CP-element group 35: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_index_resize_1/index_resize_ack
      -- CP-element group 35: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_index_scale_1/$entry
      -- CP-element group 35: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_index_scale_1/$exit
      -- CP-element group 35: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_index_scale_1/scale_rename_req
      -- CP-element group 35: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_index_scale_1/scale_rename_ack
      -- CP-element group 35: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_final_index_sum_regn_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_final_index_sum_regn_Sample/req
      -- 
    ca_3552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1521_inst_ack_1, ack => convTransposeA_CP_3268_elements(35)); -- 
    req_3577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(35), ack => array_obj_ref_1527_index_offset_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	52 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_final_index_sum_regn_sample_complete
      -- CP-element group 36: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_final_index_sum_regn_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_final_index_sum_regn_Sample/ack
      -- 
    ack_3578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1527_index_offset_ack_0, ack => convTransposeA_CP_3268_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	88 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (11) 
      -- CP-element group 37: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_offset_calculated
      -- CP-element group 37: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1528_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_final_index_sum_regn_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_final_index_sum_regn_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_base_plus_offset/sum_rename_req
      -- CP-element group 37: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1528_request/$entry
      -- CP-element group 37: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1528_request/req
      -- 
    ack_3583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1527_index_offset_ack_1, ack => convTransposeA_CP_3268_elements(37)); -- 
    req_3592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(37), ack => addr_of_1528_final_reg_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1528_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1528_request/$exit
      -- CP-element group 38: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1528_request/ack
      -- 
    ack_3593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1528_final_reg_ack_0, ack => convTransposeA_CP_3268_elements(38)); -- 
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	88 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (24) 
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1528_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1528_complete/$exit
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1528_complete/ack
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_base_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_word_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_base_address_resized
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_base_addr_resize/$entry
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_base_addr_resize/$exit
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_base_addr_resize/base_resize_req
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_base_addr_resize/base_resize_ack
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_word_addrgen/$entry
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_word_addrgen/$exit
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_word_addrgen/root_register_req
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_word_addrgen/root_register_ack
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Sample/word_access_start/$entry
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Sample/word_access_start/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Sample/word_access_start/word_0/rr
      -- 
    ack_3598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1528_final_reg_ack_1, ack => convTransposeA_CP_3268_elements(39)); -- 
    rr_3631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(39), ack => ptr_deref_1532_load_0_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Sample/word_access_start/$exit
      -- CP-element group 40: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Sample/word_access_start/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Sample/word_access_start/word_0/ra
      -- 
    ra_3632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1532_load_0_ack_0, ack => convTransposeA_CP_3268_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	88 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	49 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Update/word_access_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Update/word_access_complete/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Update/word_access_complete/word_0/ca
      -- CP-element group 41: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Update/ptr_deref_1532_Merge/$entry
      -- CP-element group 41: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Update/ptr_deref_1532_Merge/$exit
      -- CP-element group 41: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Update/ptr_deref_1532_Merge/merge_req
      -- CP-element group 41: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Update/ptr_deref_1532_Merge/merge_ack
      -- 
    ca_3643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1532_load_0_ack_1, ack => convTransposeA_CP_3268_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	29 
    -- CP-element group 42: 	31 
    -- CP-element group 42: 	33 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1542_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1542_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1542_Sample/rr
      -- 
    rr_3656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(42), ack => type_cast_1542_inst_req_0); -- 
    convTransposeA_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3268_elements(29) & convTransposeA_CP_3268_elements(31) & convTransposeA_CP_3268_elements(33);
      gj_convTransposeA_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3268_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1542_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1542_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1542_Sample/ra
      -- 
    ra_3657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1542_inst_ack_0, ack => convTransposeA_CP_3268_elements(43)); -- 
    -- CP-element group 44:  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	88 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (16) 
      -- CP-element group 44: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1542_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1542_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1542_Update/ca
      -- CP-element group 44: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_index_resized_1
      -- CP-element group 44: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_index_scaled_1
      -- CP-element group 44: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_index_computed_1
      -- CP-element group 44: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_index_resize_1/$entry
      -- CP-element group 44: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_index_resize_1/$exit
      -- CP-element group 44: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_index_resize_1/index_resize_req
      -- CP-element group 44: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_index_resize_1/index_resize_ack
      -- CP-element group 44: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_index_scale_1/$entry
      -- CP-element group 44: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_index_scale_1/$exit
      -- CP-element group 44: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_index_scale_1/scale_rename_req
      -- CP-element group 44: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_index_scale_1/scale_rename_ack
      -- CP-element group 44: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_final_index_sum_regn_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_final_index_sum_regn_Sample/req
      -- 
    ca_3662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1542_inst_ack_1, ack => convTransposeA_CP_3268_elements(44)); -- 
    req_3687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(44), ack => array_obj_ref_1548_index_offset_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	52 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_final_index_sum_regn_sample_complete
      -- CP-element group 45: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_final_index_sum_regn_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_final_index_sum_regn_Sample/ack
      -- 
    ack_3688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1548_index_offset_ack_0, ack => convTransposeA_CP_3268_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	88 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (11) 
      -- CP-element group 46: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1549_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_root_address_calculated
      -- CP-element group 46: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_offset_calculated
      -- CP-element group 46: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_final_index_sum_regn_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_final_index_sum_regn_Update/ack
      -- CP-element group 46: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_base_plus_offset/$entry
      -- CP-element group 46: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_base_plus_offset/$exit
      -- CP-element group 46: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_base_plus_offset/sum_rename_req
      -- CP-element group 46: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_base_plus_offset/sum_rename_ack
      -- CP-element group 46: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1549_request/$entry
      -- CP-element group 46: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1549_request/req
      -- 
    ack_3693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1548_index_offset_ack_1, ack => convTransposeA_CP_3268_elements(46)); -- 
    req_3702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(46), ack => addr_of_1549_final_reg_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1549_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1549_request/$exit
      -- CP-element group 47: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1549_request/ack
      -- 
    ack_3703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1549_final_reg_ack_0, ack => convTransposeA_CP_3268_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	88 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (19) 
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1549_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1549_complete/$exit
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1549_complete/ack
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_base_address_calculated
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_word_address_calculated
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_root_address_calculated
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_base_address_resized
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_base_addr_resize/$entry
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_base_addr_resize/$exit
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_base_addr_resize/base_resize_req
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_base_addr_resize/base_resize_ack
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_base_plus_offset/$entry
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_base_plus_offset/$exit
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_base_plus_offset/sum_rename_req
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_base_plus_offset/sum_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_word_addrgen/$entry
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_word_addrgen/$exit
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_word_addrgen/root_register_req
      -- CP-element group 48: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_word_addrgen/root_register_ack
      -- 
    ack_3708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1549_final_reg_ack_1, ack => convTransposeA_CP_3268_elements(48)); -- 
    -- CP-element group 49:  join  transition  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	41 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (9) 
      -- CP-element group 49: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Sample/ptr_deref_1552_Split/$entry
      -- CP-element group 49: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Sample/ptr_deref_1552_Split/$exit
      -- CP-element group 49: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Sample/ptr_deref_1552_Split/split_req
      -- CP-element group 49: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Sample/ptr_deref_1552_Split/split_ack
      -- CP-element group 49: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Sample/word_access_start/$entry
      -- CP-element group 49: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Sample/word_access_start/word_0/$entry
      -- CP-element group 49: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Sample/word_access_start/word_0/rr
      -- 
    rr_3746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(49), ack => ptr_deref_1552_store_0_req_0); -- 
    convTransposeA_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3268_elements(41) & convTransposeA_CP_3268_elements(48);
      gj_convTransposeA_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3268_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Sample/$exit
      -- CP-element group 50: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Sample/word_access_start/$exit
      -- CP-element group 50: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Sample/word_access_start/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Sample/word_access_start/word_0/ra
      -- 
    ra_3747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1552_store_0_ack_0, ack => convTransposeA_CP_3268_elements(50)); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	88 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Update/word_access_complete/$exit
      -- CP-element group 51: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Update/word_access_complete/word_0/$exit
      -- CP-element group 51: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Update/word_access_complete/word_0/ca
      -- 
    ca_3758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1552_store_0_ack_1, ack => convTransposeA_CP_3268_elements(51)); -- 
    -- CP-element group 52:  branch  join  transition  place  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	36 
    -- CP-element group 52: 	45 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (10) 
      -- CP-element group 52: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/$exit
      -- CP-element group 52: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565__exit__
      -- CP-element group 52: 	 branch_block_stmt_1301/if_stmt_1566__entry__
      -- CP-element group 52: 	 branch_block_stmt_1301/if_stmt_1566_dead_link/$entry
      -- CP-element group 52: 	 branch_block_stmt_1301/if_stmt_1566_eval_test/$entry
      -- CP-element group 52: 	 branch_block_stmt_1301/if_stmt_1566_eval_test/$exit
      -- CP-element group 52: 	 branch_block_stmt_1301/if_stmt_1566_eval_test/branch_req
      -- CP-element group 52: 	 branch_block_stmt_1301/R_cmp_1567_place
      -- CP-element group 52: 	 branch_block_stmt_1301/if_stmt_1566_if_link/$entry
      -- CP-element group 52: 	 branch_block_stmt_1301/if_stmt_1566_else_link/$entry
      -- 
    branch_req_3766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(52), ack => if_stmt_1566_branch_req_0); -- 
    convTransposeA_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3268_elements(36) & convTransposeA_CP_3268_elements(45) & convTransposeA_CP_3268_elements(51);
      gj_convTransposeA_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3268_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	97 
    -- CP-element group 53: 	98 
    -- CP-element group 53: 	100 
    -- CP-element group 53: 	101 
    -- CP-element group 53: 	103 
    -- CP-element group 53: 	104 
    -- CP-element group 53:  members (40) 
      -- CP-element group 53: 	 branch_block_stmt_1301/assign_stmt_1578__entry__
      -- CP-element group 53: 	 branch_block_stmt_1301/merge_stmt_1572__exit__
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1641/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/assign_stmt_1578__exit__
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1638/SplitProtocol/Sample/rr
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1638/SplitProtocol/Update/cr
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1638/SplitProtocol/Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1638/SplitProtocol/Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1638/SplitProtocol/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1638/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1628/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1635/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1644/SplitProtocol/Update/cr
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/Update/cr
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1644/SplitProtocol/Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/Sample/rr
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1644/SplitProtocol/Sample/rr
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1644/SplitProtocol/Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/if_stmt_1566_if_link/$exit
      -- CP-element group 53: 	 branch_block_stmt_1301/if_stmt_1566_if_link/if_choice_transition
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1644/SplitProtocol/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/whilex_xbody_ifx_xthen
      -- CP-element group 53: 	 branch_block_stmt_1301/assign_stmt_1578/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/assign_stmt_1578/$exit
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1644/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 53: 	 branch_block_stmt_1301/merge_stmt_1572_PhiReqMerge
      -- CP-element group 53: 	 branch_block_stmt_1301/merge_stmt_1572_PhiAck/$entry
      -- CP-element group 53: 	 branch_block_stmt_1301/merge_stmt_1572_PhiAck/$exit
      -- CP-element group 53: 	 branch_block_stmt_1301/merge_stmt_1572_PhiAck/dummy
      -- 
    if_choice_transition_3771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1566_branch_ack_1, ack => convTransposeA_CP_3268_elements(53)); -- 
    rr_4125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(53), ack => type_cast_1638_inst_req_0); -- 
    cr_4130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(53), ack => type_cast_1638_inst_req_1); -- 
    cr_4153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(53), ack => type_cast_1644_inst_req_1); -- 
    cr_4107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(53), ack => type_cast_1634_inst_req_1); -- 
    rr_4102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(53), ack => type_cast_1634_inst_req_0); -- 
    rr_4148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(53), ack => type_cast_1644_inst_req_0); -- 
    -- CP-element group 54:  fork  transition  place  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	56 
    -- CP-element group 54: 	58 
    -- CP-element group 54: 	60 
    -- CP-element group 54:  members (24) 
      -- CP-element group 54: 	 branch_block_stmt_1301/merge_stmt_1580__exit__
      -- CP-element group 54: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620__entry__
      -- CP-element group 54: 	 branch_block_stmt_1301/if_stmt_1566_else_link/$exit
      -- CP-element group 54: 	 branch_block_stmt_1301/if_stmt_1566_else_link/else_choice_transition
      -- CP-element group 54: 	 branch_block_stmt_1301/whilex_xbody_ifx_xelse
      -- CP-element group 54: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/$entry
      -- CP-element group 54: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1589_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1589_update_start_
      -- CP-element group 54: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1589_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1589_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1589_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1589_Update/cr
      -- CP-element group 54: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1598_update_start_
      -- CP-element group 54: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1598_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1598_Update/cr
      -- CP-element group 54: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1614_update_start_
      -- CP-element group 54: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1614_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1614_Update/cr
      -- CP-element group 54: 	 branch_block_stmt_1301/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_1301/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 54: 	 branch_block_stmt_1301/merge_stmt_1580_PhiReqMerge
      -- CP-element group 54: 	 branch_block_stmt_1301/merge_stmt_1580_PhiAck/$entry
      -- CP-element group 54: 	 branch_block_stmt_1301/merge_stmt_1580_PhiAck/$exit
      -- CP-element group 54: 	 branch_block_stmt_1301/merge_stmt_1580_PhiAck/dummy
      -- 
    else_choice_transition_3775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1566_branch_ack_0, ack => convTransposeA_CP_3268_elements(54)); -- 
    rr_3791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(54), ack => type_cast_1589_inst_req_0); -- 
    cr_3796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(54), ack => type_cast_1589_inst_req_1); -- 
    cr_3810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(54), ack => type_cast_1598_inst_req_1); -- 
    cr_3824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(54), ack => type_cast_1614_inst_req_1); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1589_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1589_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1589_Sample/ra
      -- 
    ra_3792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1589_inst_ack_0, ack => convTransposeA_CP_3268_elements(55)); -- 
    -- CP-element group 56:  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1589_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1589_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1589_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1598_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1598_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1598_Sample/rr
      -- 
    ca_3797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1589_inst_ack_1, ack => convTransposeA_CP_3268_elements(56)); -- 
    rr_3805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(56), ack => type_cast_1598_inst_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1598_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1598_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1598_Sample/ra
      -- 
    ra_3806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1598_inst_ack_0, ack => convTransposeA_CP_3268_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	54 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1598_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1598_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1598_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1614_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1614_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1614_Sample/rr
      -- 
    ca_3811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1598_inst_ack_1, ack => convTransposeA_CP_3268_elements(58)); -- 
    rr_3819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(58), ack => type_cast_1614_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1614_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1614_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1614_Sample/ra
      -- 
    ra_3820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1614_inst_ack_0, ack => convTransposeA_CP_3268_elements(59)); -- 
    -- CP-element group 60:  branch  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	54 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (13) 
      -- CP-element group 60: 	 branch_block_stmt_1301/if_stmt_1621__entry__
      -- CP-element group 60: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620__exit__
      -- CP-element group 60: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/$exit
      -- CP-element group 60: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1614_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1614_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1301/assign_stmt_1586_to_assign_stmt_1620/type_cast_1614_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_1301/if_stmt_1621_dead_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_1301/if_stmt_1621_eval_test/$entry
      -- CP-element group 60: 	 branch_block_stmt_1301/if_stmt_1621_eval_test/$exit
      -- CP-element group 60: 	 branch_block_stmt_1301/if_stmt_1621_eval_test/branch_req
      -- CP-element group 60: 	 branch_block_stmt_1301/R_cmp111_1622_place
      -- CP-element group 60: 	 branch_block_stmt_1301/if_stmt_1621_if_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_1301/if_stmt_1621_else_link/$entry
      -- 
    ca_3825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1614_inst_ack_1, ack => convTransposeA_CP_3268_elements(60)); -- 
    branch_req_3833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(60), ack => if_stmt_1621_branch_req_0); -- 
    -- CP-element group 61:  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (15) 
      -- CP-element group 61: 	 branch_block_stmt_1301/merge_stmt_1655__exit__
      -- CP-element group 61: 	 branch_block_stmt_1301/assign_stmt_1660__entry__
      -- CP-element group 61: 	 branch_block_stmt_1301/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_1301/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 61: 	 branch_block_stmt_1301/merge_stmt_1655_PhiAck/$entry
      -- CP-element group 61: 	 branch_block_stmt_1301/merge_stmt_1655_PhiAck/$exit
      -- CP-element group 61: 	 branch_block_stmt_1301/merge_stmt_1655_PhiAck/dummy
      -- CP-element group 61: 	 branch_block_stmt_1301/merge_stmt_1655_PhiReqMerge
      -- CP-element group 61: 	 branch_block_stmt_1301/if_stmt_1621_if_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_1301/if_stmt_1621_if_link/if_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_1301/ifx_xelse_whilex_xend
      -- CP-element group 61: 	 branch_block_stmt_1301/assign_stmt_1660/$entry
      -- CP-element group 61: 	 branch_block_stmt_1301/assign_stmt_1660/WPIPE_Block0_done_1657_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_1301/assign_stmt_1660/WPIPE_Block0_done_1657_Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_1301/assign_stmt_1660/WPIPE_Block0_done_1657_Sample/req
      -- 
    if_choice_transition_3838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1621_branch_ack_1, ack => convTransposeA_CP_3268_elements(61)); -- 
    req_3858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(61), ack => WPIPE_Block0_done_1657_inst_req_0); -- 
    -- CP-element group 62:  fork  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	89 
    -- CP-element group 62: 	90 
    -- CP-element group 62: 	91 
    -- CP-element group 62: 	93 
    -- CP-element group 62: 	94 
    -- CP-element group 62:  members (22) 
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1646/SplitProtocol/Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1635/$entry
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1646/SplitProtocol/$entry
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/$entry
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1640/$entry
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1646/$entry
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/$entry
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1646/SplitProtocol/Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1640/SplitProtocol/$entry
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1640/SplitProtocol/Update/cr
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/$entry
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1641/$entry
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1646/SplitProtocol/Update/cr
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1628/$entry
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1640/SplitProtocol/Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1640/SplitProtocol/Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1640/SplitProtocol/Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1646/SplitProtocol/Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/$entry
      -- CP-element group 62: 	 branch_block_stmt_1301/if_stmt_1621_else_link/$exit
      -- CP-element group 62: 	 branch_block_stmt_1301/if_stmt_1621_else_link/else_choice_transition
      -- CP-element group 62: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122
      -- 
    else_choice_transition_3842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1621_branch_ack_0, ack => convTransposeA_CP_3268_elements(62)); -- 
    rr_4076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(62), ack => type_cast_1646_inst_req_0); -- 
    cr_4058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(62), ack => type_cast_1640_inst_req_1); -- 
    cr_4081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(62), ack => type_cast_1646_inst_req_1); -- 
    rr_4053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(62), ack => type_cast_1640_inst_req_0); -- 
    -- CP-element group 63:  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_1301/assign_stmt_1660/WPIPE_Block0_done_1657_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1301/assign_stmt_1660/WPIPE_Block0_done_1657_update_start_
      -- CP-element group 63: 	 branch_block_stmt_1301/assign_stmt_1660/WPIPE_Block0_done_1657_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1301/assign_stmt_1660/WPIPE_Block0_done_1657_Sample/ack
      -- CP-element group 63: 	 branch_block_stmt_1301/assign_stmt_1660/WPIPE_Block0_done_1657_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_1301/assign_stmt_1660/WPIPE_Block0_done_1657_Update/req
      -- 
    ack_3859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1657_inst_ack_0, ack => convTransposeA_CP_3268_elements(63)); -- 
    req_3863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(63), ack => WPIPE_Block0_done_1657_inst_req_1); -- 
    -- CP-element group 64:  transition  place  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (16) 
      -- CP-element group 64: 	 branch_block_stmt_1301/$exit
      -- CP-element group 64: 	 $exit
      -- CP-element group 64: 	 branch_block_stmt_1301/branch_block_stmt_1301__exit__
      -- CP-element group 64: 	 branch_block_stmt_1301/assign_stmt_1660__exit__
      -- CP-element group 64: 	 branch_block_stmt_1301/return__
      -- CP-element group 64: 	 branch_block_stmt_1301/merge_stmt_1662__exit__
      -- CP-element group 64: 	 branch_block_stmt_1301/merge_stmt_1662_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_1301/return___PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_1301/merge_stmt_1662_PhiAck/dummy
      -- CP-element group 64: 	 branch_block_stmt_1301/merge_stmt_1662_PhiAck/$exit
      -- CP-element group 64: 	 branch_block_stmt_1301/merge_stmt_1662_PhiAck/$entry
      -- CP-element group 64: 	 branch_block_stmt_1301/return___PhiReq/$exit
      -- CP-element group 64: 	 branch_block_stmt_1301/assign_stmt_1660/$exit
      -- CP-element group 64: 	 branch_block_stmt_1301/assign_stmt_1660/WPIPE_Block0_done_1657_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1301/assign_stmt_1660/WPIPE_Block0_done_1657_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1301/assign_stmt_1660/WPIPE_Block0_done_1657_Update/ack
      -- 
    ack_3864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1657_inst_ack_1, ack => convTransposeA_CP_3268_elements(64)); -- 
    -- CP-element group 65:  transition  output  delay-element  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	27 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	69 
    -- CP-element group 65:  members (4) 
      -- CP-element group 65: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1408/$exit
      -- CP-element group 65: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/$exit
      -- CP-element group 65: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1412_konst_delay_trans
      -- CP-element group 65: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_req
      -- 
    phi_stmt_1408_req_3875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1408_req_3875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(65), ack => phi_stmt_1408_req_0); -- 
    -- Element group convTransposeA_CP_3268_elements(65) is a control-delay.
    cp_element_65_delay: control_delay_element  generic map(name => " 65_delay", delay_value => 1)  port map(req => convTransposeA_CP_3268_elements(27), ack => convTransposeA_CP_3268_elements(65), clk => clk, reset =>reset);
    -- CP-element group 66:  transition  output  delay-element  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	27 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	69 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1415/$exit
      -- CP-element group 66: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_sources/$exit
      -- CP-element group 66: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_sources/type_cast_1420_konst_delay_trans
      -- CP-element group 66: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_req
      -- 
    phi_stmt_1415_req_3883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1415_req_3883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(66), ack => phi_stmt_1415_req_0); -- 
    -- Element group convTransposeA_CP_3268_elements(66) is a control-delay.
    cp_element_66_delay: control_delay_element  generic map(name => " 66_delay", delay_value => 1)  port map(req => convTransposeA_CP_3268_elements(27), ack => convTransposeA_CP_3268_elements(66), clk => clk, reset =>reset);
    -- CP-element group 67:  transition  output  delay-element  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	27 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1423/$exit
      -- CP-element group 67: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/$exit
      -- CP-element group 67: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1427_konst_delay_trans
      -- CP-element group 67: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_req
      -- 
    phi_stmt_1423_req_3891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1423_req_3891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(67), ack => phi_stmt_1423_req_0); -- 
    -- Element group convTransposeA_CP_3268_elements(67) is a control-delay.
    cp_element_67_delay: control_delay_element  generic map(name => " 67_delay", delay_value => 1)  port map(req => convTransposeA_CP_3268_elements(27), ack => convTransposeA_CP_3268_elements(67), clk => clk, reset =>reset);
    -- CP-element group 68:  transition  output  delay-element  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	27 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1430/$exit
      -- CP-element group 68: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_sources/$exit
      -- CP-element group 68: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_sources/type_cast_1434_konst_delay_trans
      -- CP-element group 68: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_req
      -- 
    phi_stmt_1430_req_3899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1430_req_3899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(68), ack => phi_stmt_1430_req_0); -- 
    -- Element group convTransposeA_CP_3268_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => convTransposeA_CP_3268_elements(27), ack => convTransposeA_CP_3268_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  join  transition  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	65 
    -- CP-element group 69: 	66 
    -- CP-element group 69: 	67 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	83 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1301/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3268_elements(65) & convTransposeA_CP_3268_elements(66) & convTransposeA_CP_3268_elements(67) & convTransposeA_CP_3268_elements(68);
      gj_convTransposeA_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3268_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	1 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1414/SplitProtocol/Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1414/SplitProtocol/Sample/ra
      -- 
    ra_3919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1414_inst_ack_0, ack => convTransposeA_CP_3268_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	1 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1414/SplitProtocol/Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1414/SplitProtocol/Update/ca
      -- 
    ca_3924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1414_inst_ack_1, ack => convTransposeA_CP_3268_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	82 
    -- CP-element group 72:  members (5) 
      -- CP-element group 72: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1408/$exit
      -- CP-element group 72: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/$exit
      -- CP-element group 72: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1414/$exit
      -- CP-element group 72: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_sources/type_cast_1414/SplitProtocol/$exit
      -- CP-element group 72: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1408/phi_stmt_1408_req
      -- 
    phi_stmt_1408_req_3925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1408_req_3925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(72), ack => phi_stmt_1408_req_1); -- 
    convTransposeA_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3268_elements(70) & convTransposeA_CP_3268_elements(71);
      gj_convTransposeA_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3268_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	1 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_sources/type_cast_1422/SplitProtocol/Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_sources/type_cast_1422/SplitProtocol/Sample/ra
      -- 
    ra_3942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1422_inst_ack_0, ack => convTransposeA_CP_3268_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	1 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_sources/type_cast_1422/SplitProtocol/Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_sources/type_cast_1422/SplitProtocol/Update/ca
      -- 
    ca_3947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1422_inst_ack_1, ack => convTransposeA_CP_3268_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	82 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1415/$exit
      -- CP-element group 75: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_sources/$exit
      -- CP-element group 75: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_sources/type_cast_1422/$exit
      -- CP-element group 75: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_sources/type_cast_1422/SplitProtocol/$exit
      -- CP-element group 75: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1415/phi_stmt_1415_req
      -- 
    phi_stmt_1415_req_3948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1415_req_3948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(75), ack => phi_stmt_1415_req_1); -- 
    convTransposeA_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3268_elements(73) & convTransposeA_CP_3268_elements(74);
      gj_convTransposeA_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3268_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	1 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Sample/ra
      -- 
    ra_3965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1429_inst_ack_0, ack => convTransposeA_CP_3268_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	1 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/Update/ca
      -- 
    ca_3970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1429_inst_ack_1, ack => convTransposeA_CP_3268_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	82 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1423/$exit
      -- CP-element group 78: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/$exit
      -- CP-element group 78: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/$exit
      -- CP-element group 78: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_sources/type_cast_1429/SplitProtocol/$exit
      -- CP-element group 78: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1423/phi_stmt_1423_req
      -- 
    phi_stmt_1423_req_3971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1423_req_3971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(78), ack => phi_stmt_1423_req_1); -- 
    convTransposeA_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3268_elements(76) & convTransposeA_CP_3268_elements(77);
      gj_convTransposeA_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3268_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	1 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_sources/type_cast_1436/SplitProtocol/Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_sources/type_cast_1436/SplitProtocol/Sample/ra
      -- 
    ra_3988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1436_inst_ack_0, ack => convTransposeA_CP_3268_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	1 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_sources/type_cast_1436/SplitProtocol/Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_sources/type_cast_1436/SplitProtocol/Update/ca
      -- 
    ca_3993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1436_inst_ack_1, ack => convTransposeA_CP_3268_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1430/$exit
      -- CP-element group 81: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_sources/type_cast_1436/$exit
      -- CP-element group 81: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_sources/type_cast_1436/SplitProtocol/$exit
      -- CP-element group 81: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/phi_stmt_1430/phi_stmt_1430_req
      -- 
    phi_stmt_1430_req_3994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1430_req_3994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(81), ack => phi_stmt_1430_req_1); -- 
    convTransposeA_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3268_elements(79) & convTransposeA_CP_3268_elements(80);
      gj_convTransposeA_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3268_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  join  transition  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	72 
    -- CP-element group 82: 	75 
    -- CP-element group 82: 	78 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1301/ifx_xend122_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3268_elements(72) & convTransposeA_CP_3268_elements(75) & convTransposeA_CP_3268_elements(78) & convTransposeA_CP_3268_elements(81);
      gj_convTransposeA_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3268_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  merge  fork  transition  place  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	69 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	85 
    -- CP-element group 83: 	86 
    -- CP-element group 83: 	87 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1301/merge_stmt_1407_PhiReqMerge
      -- CP-element group 83: 	 branch_block_stmt_1301/merge_stmt_1407_PhiAck/$entry
      -- 
    convTransposeA_CP_3268_elements(83) <= OrReduce(convTransposeA_CP_3268_elements(69) & convTransposeA_CP_3268_elements(82));
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	88 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1301/merge_stmt_1407_PhiAck/phi_stmt_1408_ack
      -- 
    phi_stmt_1408_ack_3999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1408_ack_0, ack => convTransposeA_CP_3268_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	88 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1301/merge_stmt_1407_PhiAck/phi_stmt_1415_ack
      -- 
    phi_stmt_1415_ack_4000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1415_ack_0, ack => convTransposeA_CP_3268_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_1301/merge_stmt_1407_PhiAck/phi_stmt_1423_ack
      -- 
    phi_stmt_1423_ack_4001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1423_ack_0, ack => convTransposeA_CP_3268_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	83 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_1301/merge_stmt_1407_PhiAck/phi_stmt_1430_ack
      -- 
    phi_stmt_1430_ack_4002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1430_ack_0, ack => convTransposeA_CP_3268_elements(87)); -- 
    -- CP-element group 88:  join  fork  transition  place  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	84 
    -- CP-element group 88: 	85 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	28 
    -- CP-element group 88: 	29 
    -- CP-element group 88: 	30 
    -- CP-element group 88: 	31 
    -- CP-element group 88: 	32 
    -- CP-element group 88: 	33 
    -- CP-element group 88: 	34 
    -- CP-element group 88: 	35 
    -- CP-element group 88: 	37 
    -- CP-element group 88: 	39 
    -- CP-element group 88: 	41 
    -- CP-element group 88: 	44 
    -- CP-element group 88: 	46 
    -- CP-element group 88: 	48 
    -- CP-element group 88: 	51 
    -- CP-element group 88:  members (53) 
      -- CP-element group 88: 	 branch_block_stmt_1301/merge_stmt_1407__exit__
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1451_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1451_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1465_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1465_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565__entry__
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1465_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1465_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1465_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1451_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1521_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1479_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1479_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1451_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1479_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1521_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1521_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1521_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1521_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1451_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1528_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1479_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1465_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1521_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1479_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1479_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1451_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_final_index_sum_regn_update_start
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_final_index_sum_regn_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1527_final_index_sum_regn_Update/req
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1528_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1528_complete/req
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Update/word_access_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Update/word_access_complete/word_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1532_Update/word_access_complete/word_0/cr
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1542_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1542_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/type_cast_1542_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1549_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_final_index_sum_regn_update_start
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_final_index_sum_regn_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/array_obj_ref_1548_final_index_sum_regn_Update/req
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1549_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/addr_of_1549_complete/req
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Update/word_access_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Update/word_access_complete/word_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_1301/assign_stmt_1443_to_assign_stmt_1565/ptr_deref_1552_Update/word_access_complete/word_0/cr
      -- CP-element group 88: 	 branch_block_stmt_1301/merge_stmt_1407_PhiAck/$exit
      -- 
    cr_3523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(88), ack => type_cast_1465_inst_req_1); -- 
    rr_3518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(88), ack => type_cast_1465_inst_req_0); -- 
    cr_3551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(88), ack => type_cast_1521_inst_req_1); -- 
    rr_3532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(88), ack => type_cast_1479_inst_req_0); -- 
    cr_3509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(88), ack => type_cast_1451_inst_req_1); -- 
    cr_3537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(88), ack => type_cast_1479_inst_req_1); -- 
    rr_3546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(88), ack => type_cast_1521_inst_req_0); -- 
    rr_3504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(88), ack => type_cast_1451_inst_req_0); -- 
    req_3582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(88), ack => array_obj_ref_1527_index_offset_req_1); -- 
    req_3597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(88), ack => addr_of_1528_final_reg_req_1); -- 
    cr_3642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(88), ack => ptr_deref_1532_load_0_req_1); -- 
    cr_3661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(88), ack => type_cast_1542_inst_req_1); -- 
    req_3692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(88), ack => array_obj_ref_1548_index_offset_req_1); -- 
    req_3707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(88), ack => addr_of_1549_final_reg_req_1); -- 
    cr_3757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(88), ack => ptr_deref_1552_store_0_req_1); -- 
    convTransposeA_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3268_elements(84) & convTransposeA_CP_3268_elements(85) & convTransposeA_CP_3268_elements(86) & convTransposeA_CP_3268_elements(87);
      gj_convTransposeA_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3268_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  output  delay-element  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	62 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	96 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_req
      -- CP-element group 89: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1632_konst_delay_trans
      -- CP-element group 89: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1628/$exit
      -- 
    phi_stmt_1628_req_4037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1628_req_4037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(89), ack => phi_stmt_1628_req_0); -- 
    -- Element group convTransposeA_CP_3268_elements(89) is a control-delay.
    cp_element_89_delay: control_delay_element  generic map(name => " 89_delay", delay_value => 1)  port map(req => convTransposeA_CP_3268_elements(62), ack => convTransposeA_CP_3268_elements(89), clk => clk, reset =>reset);
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	62 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1640/SplitProtocol/Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1640/SplitProtocol/Sample/$exit
      -- 
    ra_4054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1640_inst_ack_0, ack => convTransposeA_CP_3268_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	62 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1640/SplitProtocol/Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1640/SplitProtocol/Update/ca
      -- 
    ca_4059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1640_inst_ack_1, ack => convTransposeA_CP_3268_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	96 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1635/$exit
      -- CP-element group 92: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1640/$exit
      -- CP-element group 92: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_req
      -- CP-element group 92: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1640/SplitProtocol/$exit
      -- 
    phi_stmt_1635_req_4060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1635_req_4060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(92), ack => phi_stmt_1635_req_1); -- 
    convTransposeA_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3268_elements(90) & convTransposeA_CP_3268_elements(91);
      gj_convTransposeA_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3268_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	62 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1646/SplitProtocol/Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1646/SplitProtocol/Sample/ra
      -- 
    ra_4077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1646_inst_ack_0, ack => convTransposeA_CP_3268_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	62 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1646/SplitProtocol/Update/ca
      -- CP-element group 94: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1646/SplitProtocol/Update/$exit
      -- 
    ca_4082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1646_inst_ack_1, ack => convTransposeA_CP_3268_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1646/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1646/$exit
      -- CP-element group 95: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1641/$exit
      -- CP-element group 95: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_req
      -- 
    phi_stmt_1641_req_4083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1641_req_4083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(95), ack => phi_stmt_1641_req_1); -- 
    convTransposeA_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3268_elements(93) & convTransposeA_CP_3268_elements(94);
      gj_convTransposeA_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3268_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	89 
    -- CP-element group 96: 	92 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	107 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_1301/ifx_xelse_ifx_xend122_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3268_elements(89) & convTransposeA_CP_3268_elements(92) & convTransposeA_CP_3268_elements(95);
      gj_convTransposeA_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3268_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	53 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/Sample/ra
      -- CP-element group 97: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/Sample/$exit
      -- 
    ra_4103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1634_inst_ack_0, ack => convTransposeA_CP_3268_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	53 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/Update/ca
      -- CP-element group 98: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/Update/$exit
      -- 
    ca_4108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1634_inst_ack_1, ack => convTransposeA_CP_3268_elements(98)); -- 
    -- CP-element group 99:  join  transition  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	106 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/$exit
      -- CP-element group 99: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1628/$exit
      -- CP-element group 99: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_req
      -- CP-element group 99: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/SplitProtocol/$exit
      -- CP-element group 99: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1628/phi_stmt_1628_sources/type_cast_1634/$exit
      -- 
    phi_stmt_1628_req_4109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1628_req_4109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(99), ack => phi_stmt_1628_req_1); -- 
    convTransposeA_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3268_elements(97) & convTransposeA_CP_3268_elements(98);
      gj_convTransposeA_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3268_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	53 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1638/SplitProtocol/Sample/ra
      -- CP-element group 100: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1638/SplitProtocol/Sample/$exit
      -- 
    ra_4126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1638_inst_ack_0, ack => convTransposeA_CP_3268_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	53 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1638/SplitProtocol/Update/ca
      -- CP-element group 101: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1638/SplitProtocol/Update/$exit
      -- 
    ca_4131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1638_inst_ack_1, ack => convTransposeA_CP_3268_elements(101)); -- 
    -- CP-element group 102:  join  transition  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	106 
    -- CP-element group 102:  members (5) 
      -- CP-element group 102: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_req
      -- CP-element group 102: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1638/SplitProtocol/$exit
      -- CP-element group 102: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/type_cast_1638/$exit
      -- CP-element group 102: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1635/phi_stmt_1635_sources/$exit
      -- CP-element group 102: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1635/$exit
      -- 
    phi_stmt_1635_req_4132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1635_req_4132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(102), ack => phi_stmt_1635_req_0); -- 
    convTransposeA_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3268_elements(100) & convTransposeA_CP_3268_elements(101);
      gj_convTransposeA_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3268_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	53 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1644/SplitProtocol/Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1644/SplitProtocol/Sample/$exit
      -- 
    ra_4149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1644_inst_ack_0, ack => convTransposeA_CP_3268_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	53 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1644/SplitProtocol/Update/ca
      -- CP-element group 104: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1644/SplitProtocol/Update/$exit
      -- 
    ca_4154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1644_inst_ack_1, ack => convTransposeA_CP_3268_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (5) 
      -- CP-element group 105: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1641/$exit
      -- CP-element group 105: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_req
      -- CP-element group 105: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1644/SplitProtocol/$exit
      -- CP-element group 105: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/type_cast_1644/$exit
      -- CP-element group 105: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/phi_stmt_1641/phi_stmt_1641_sources/$exit
      -- 
    phi_stmt_1641_req_4155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1641_req_4155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3268_elements(105), ack => phi_stmt_1641_req_0); -- 
    convTransposeA_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3268_elements(103) & convTransposeA_CP_3268_elements(104);
      gj_convTransposeA_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3268_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  join  transition  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	99 
    -- CP-element group 106: 	102 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_1301/ifx_xthen_ifx_xend122_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3268_elements(99) & convTransposeA_CP_3268_elements(102) & convTransposeA_CP_3268_elements(105);
      gj_convTransposeA_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3268_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  merge  fork  transition  place  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	96 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	109 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1301/merge_stmt_1627_PhiAck/$entry
      -- CP-element group 107: 	 branch_block_stmt_1301/merge_stmt_1627_PhiReqMerge
      -- 
    convTransposeA_CP_3268_elements(107) <= OrReduce(convTransposeA_CP_3268_elements(96) & convTransposeA_CP_3268_elements(106));
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	111 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_1301/merge_stmt_1627_PhiAck/phi_stmt_1628_ack
      -- 
    phi_stmt_1628_ack_4160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1628_ack_0, ack => convTransposeA_CP_3268_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_1301/merge_stmt_1627_PhiAck/phi_stmt_1635_ack
      -- 
    phi_stmt_1635_ack_4161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1635_ack_0, ack => convTransposeA_CP_3268_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1301/merge_stmt_1627_PhiAck/phi_stmt_1641_ack
      -- 
    phi_stmt_1641_ack_4162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1641_ack_0, ack => convTransposeA_CP_3268_elements(110)); -- 
    -- CP-element group 111:  join  transition  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	108 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	1 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_1301/merge_stmt_1627_PhiAck/$exit
      -- 
    convTransposeA_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeA_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeA_CP_3268_elements(108) & convTransposeA_CP_3268_elements(109) & convTransposeA_CP_3268_elements(110);
      gj_convTransposeA_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3268_elements(111), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom80_1547_resized : std_logic_vector(13 downto 0);
    signal R_idxprom80_1547_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1526_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1526_scaled : std_logic_vector(13 downto 0);
    signal add53_1364 : std_logic_vector(31 downto 0);
    signal add72_1502 : std_logic_vector(31 downto 0);
    signal add74_1512 : std_logic_vector(31 downto 0);
    signal add85_1560 : std_logic_vector(31 downto 0);
    signal add92_1578 : std_logic_vector(15 downto 0);
    signal add_1353 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_1448 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1527_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1527_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1527_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1527_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1527_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1527_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1548_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1548_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1548_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1548_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1548_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1548_root_address : std_logic_vector(13 downto 0);
    signal arrayidx76_1529 : std_logic_vector(31 downto 0);
    signal arrayidx81_1550 : std_logic_vector(31 downto 0);
    signal call10_1316 : std_logic_vector(31 downto 0);
    signal call13_1319 : std_logic_vector(31 downto 0);
    signal call16_1322 : std_logic_vector(31 downto 0);
    signal call19_1325 : std_logic_vector(31 downto 0);
    signal call1_1307 : std_logic_vector(31 downto 0);
    signal call21_1328 : std_logic_vector(31 downto 0);
    signal call23_1331 : std_logic_vector(31 downto 0);
    signal call24_1334 : std_logic_vector(31 downto 0);
    signal call27_1337 : std_logic_vector(31 downto 0);
    signal call30_1340 : std_logic_vector(31 downto 0);
    signal call4_1310 : std_logic_vector(31 downto 0);
    signal call7_1313 : std_logic_vector(31 downto 0);
    signal call_1304 : std_logic_vector(31 downto 0);
    signal cmp100_1595 : std_logic_vector(0 downto 0);
    signal cmp111_1620 : std_logic_vector(0 downto 0);
    signal cmp_1565 : std_logic_vector(0 downto 0);
    signal conv106_1615 : std_logic_vector(31 downto 0);
    signal conv109_1399 : std_logic_vector(31 downto 0);
    signal conv35_1452 : std_logic_vector(31 downto 0);
    signal conv37_1347 : std_logic_vector(31 downto 0);
    signal conv46_1466 : std_logic_vector(31 downto 0);
    signal conv60_1480 : std_logic_vector(31 downto 0);
    signal conv63_1375 : std_logic_vector(31 downto 0);
    signal conv65_1486 : std_logic_vector(31 downto 0);
    signal conv68_1381 : std_logic_vector(31 downto 0);
    signal conv70_1492 : std_logic_vector(31 downto 0);
    signal conv88_1387 : std_logic_vector(31 downto 0);
    signal conv96_1590 : std_logic_vector(31 downto 0);
    signal conv99_1393 : std_logic_vector(31 downto 0);
    signal idxprom80_1543 : std_logic_vector(63 downto 0);
    signal idxprom_1522 : std_logic_vector(63 downto 0);
    signal inc104_1599 : std_logic_vector(15 downto 0);
    signal inc104x_xinput_dim0x_x2_1604 : std_logic_vector(15 downto 0);
    signal inc_1586 : std_logic_vector(15 downto 0);
    signal indvar_1408 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_1653 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_1641 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1430 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_1635 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1423 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1611 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_1628 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1415 : std_logic_vector(15 downto 0);
    signal mul49_1471 : std_logic_vector(31 downto 0);
    signal mul71_1497 : std_logic_vector(31 downto 0);
    signal mul73_1507 : std_logic_vector(31 downto 0);
    signal mul_1457 : std_logic_vector(31 downto 0);
    signal ptr_deref_1532_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1532_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1532_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1532_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1532_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1552_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1552_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1552_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1552_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1552_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1552_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr110125_1405 : std_logic_vector(31 downto 0);
    signal shr79_1539 : std_logic_vector(31 downto 0);
    signal shr_1518 : std_logic_vector(31 downto 0);
    signal sub43_1462 : std_logic_vector(31 downto 0);
    signal sub56_1369 : std_logic_vector(31 downto 0);
    signal sub57_1476 : std_logic_vector(31 downto 0);
    signal sub_1358 : std_logic_vector(31 downto 0);
    signal tmp1_1443 : std_logic_vector(31 downto 0);
    signal tmp77_1533 : std_logic_vector(63 downto 0);
    signal type_cast_1345_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1351_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1362_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1373_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1379_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1385_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1391_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1397_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1403_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1412_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1414_wire : std_logic_vector(31 downto 0);
    signal type_cast_1420_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1422_wire : std_logic_vector(15 downto 0);
    signal type_cast_1427_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1429_wire : std_logic_vector(15 downto 0);
    signal type_cast_1434_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1436_wire : std_logic_vector(15 downto 0);
    signal type_cast_1441_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1484_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1490_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1516_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1537_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1558_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1576_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1584_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1608_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1632_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1634_wire : std_logic_vector(15 downto 0);
    signal type_cast_1638_wire : std_logic_vector(15 downto 0);
    signal type_cast_1640_wire : std_logic_vector(15 downto 0);
    signal type_cast_1644_wire : std_logic_vector(15 downto 0);
    signal type_cast_1646_wire : std_logic_vector(15 downto 0);
    signal type_cast_1651_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1659_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1527_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1527_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1527_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1527_resized_base_address <= "00000000000000";
    array_obj_ref_1548_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1548_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1548_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1548_resized_base_address <= "00000000000000";
    ptr_deref_1532_word_offset_0 <= "00000000000000";
    ptr_deref_1552_word_offset_0 <= "00000000000000";
    type_cast_1345_wire_constant <= "00000000000000001111111111111111";
    type_cast_1351_wire_constant <= "00000000000000001111111111111111";
    type_cast_1362_wire_constant <= "00000000000000001111111111111111";
    type_cast_1373_wire_constant <= "00000000000000001111111111111111";
    type_cast_1379_wire_constant <= "00000000000000001111111111111111";
    type_cast_1385_wire_constant <= "00000000000000001111111111111111";
    type_cast_1391_wire_constant <= "00000000000000001111111111111111";
    type_cast_1397_wire_constant <= "00000000000000000000000000000010";
    type_cast_1403_wire_constant <= "00000000000000000011111111111111";
    type_cast_1412_wire_constant <= "00000000000000000000000000000000";
    type_cast_1420_wire_constant <= "0000000000000000";
    type_cast_1427_wire_constant <= "0000000000000000";
    type_cast_1434_wire_constant <= "0000000000000000";
    type_cast_1441_wire_constant <= "00000000000000000000000000000100";
    type_cast_1484_wire_constant <= "00000000000000001111111111111111";
    type_cast_1490_wire_constant <= "00000000000000001111111111111111";
    type_cast_1516_wire_constant <= "00000000000000000000000000000010";
    type_cast_1537_wire_constant <= "00000000000000000000000000000010";
    type_cast_1558_wire_constant <= "00000000000000000000000000000100";
    type_cast_1576_wire_constant <= "0000000000000100";
    type_cast_1584_wire_constant <= "0000000000000001";
    type_cast_1608_wire_constant <= "0000000000000000";
    type_cast_1632_wire_constant <= "0000000000000000";
    type_cast_1651_wire_constant <= "00000000000000000000000000000001";
    type_cast_1659_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_1408: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1412_wire_constant & type_cast_1414_wire;
      req <= phi_stmt_1408_req_0 & phi_stmt_1408_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1408",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1408_ack_0,
          idata => idata,
          odata => indvar_1408,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1408
    phi_stmt_1415: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1420_wire_constant & type_cast_1422_wire;
      req <= phi_stmt_1415_req_0 & phi_stmt_1415_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1415",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1415_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1415,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1415
    phi_stmt_1423: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1427_wire_constant & type_cast_1429_wire;
      req <= phi_stmt_1423_req_0 & phi_stmt_1423_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1423",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1423_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1423,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1423
    phi_stmt_1430: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1434_wire_constant & type_cast_1436_wire;
      req <= phi_stmt_1430_req_0 & phi_stmt_1430_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1430",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1430_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1430,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1430
    phi_stmt_1628: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1632_wire_constant & type_cast_1634_wire;
      req <= phi_stmt_1628_req_0 & phi_stmt_1628_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1628",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1628_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_1628,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1628
    phi_stmt_1635: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1638_wire & type_cast_1640_wire;
      req <= phi_stmt_1635_req_0 & phi_stmt_1635_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1635",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1635_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_1635,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1635
    phi_stmt_1641: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1644_wire & type_cast_1646_wire;
      req <= phi_stmt_1641_req_0 & phi_stmt_1641_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1641",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1641_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_1641,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1641
    -- flow-through select operator MUX_1610_inst
    input_dim1x_x2_1611 <= type_cast_1608_wire_constant when (cmp100_1595(0) /=  '0') else inc_1586;
    addr_of_1528_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1528_final_reg_req_0;
      addr_of_1528_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1528_final_reg_req_1;
      addr_of_1528_final_reg_ack_1<= rack(0);
      addr_of_1528_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1528_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1527_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx76_1529,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1549_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1549_final_reg_req_0;
      addr_of_1549_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1549_final_reg_req_1;
      addr_of_1549_final_reg_ack_1<= rack(0);
      addr_of_1549_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1549_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1548_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx81_1550,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1414_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1414_inst_req_0;
      type_cast_1414_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1414_inst_req_1;
      type_cast_1414_inst_ack_1<= rack(0);
      type_cast_1414_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1414_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1653,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1414_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1422_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1422_inst_req_0;
      type_cast_1422_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1422_inst_req_1;
      type_cast_1422_inst_ack_1<= rack(0);
      type_cast_1422_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1422_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_1628,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1422_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1429_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1429_inst_req_0;
      type_cast_1429_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1429_inst_req_1;
      type_cast_1429_inst_ack_1<= rack(0);
      type_cast_1429_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1429_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_1635,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1429_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1436_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1436_inst_req_0;
      type_cast_1436_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1436_inst_req_1;
      type_cast_1436_inst_ack_1<= rack(0);
      type_cast_1436_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1436_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_1641,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1436_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1451_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1451_inst_req_0;
      type_cast_1451_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1451_inst_req_1;
      type_cast_1451_inst_ack_1<= rack(0);
      type_cast_1451_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1451_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1430,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_1452,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1465_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1465_inst_req_0;
      type_cast_1465_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1465_inst_req_1;
      type_cast_1465_inst_ack_1<= rack(0);
      type_cast_1465_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1465_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1423,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv46_1466,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1479_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1479_inst_req_0;
      type_cast_1479_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1479_inst_req_1;
      type_cast_1479_inst_ack_1<= rack(0);
      type_cast_1479_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1479_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1415,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv60_1480,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1521_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1521_inst_req_0;
      type_cast_1521_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1521_inst_req_1;
      type_cast_1521_inst_ack_1<= rack(0);
      type_cast_1521_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1521_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr_1518,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1522,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1542_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1542_inst_req_0;
      type_cast_1542_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1542_inst_req_1;
      type_cast_1542_inst_ack_1<= rack(0);
      type_cast_1542_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1542_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr79_1539,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom80_1543,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1589_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1589_inst_req_0;
      type_cast_1589_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1589_inst_req_1;
      type_cast_1589_inst_ack_1<= rack(0);
      type_cast_1589_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1589_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_1586,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv96_1590,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1598_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1598_inst_req_0;
      type_cast_1598_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1598_inst_req_1;
      type_cast_1598_inst_ack_1<= rack(0);
      type_cast_1598_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1598_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp100_1595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc104_1599,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1614_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1614_inst_req_0;
      type_cast_1614_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1614_inst_req_1;
      type_cast_1614_inst_ack_1<= rack(0);
      type_cast_1614_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1614_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc104x_xinput_dim0x_x2_1604,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv106_1615,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1634_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1634_inst_req_0;
      type_cast_1634_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1634_inst_req_1;
      type_cast_1634_inst_ack_1<= rack(0);
      type_cast_1634_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1634_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add92_1578,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1634_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1638_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1638_inst_req_0;
      type_cast_1638_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1638_inst_req_1;
      type_cast_1638_inst_ack_1<= rack(0);
      type_cast_1638_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1638_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1423,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1638_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1640_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1640_inst_req_0;
      type_cast_1640_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1640_inst_req_1;
      type_cast_1640_inst_ack_1<= rack(0);
      type_cast_1640_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1640_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1611,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1640_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1644_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1644_inst_req_0;
      type_cast_1644_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1644_inst_req_1;
      type_cast_1644_inst_ack_1<= rack(0);
      type_cast_1644_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1644_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1430,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1644_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1646_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1646_inst_req_0;
      type_cast_1646_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1646_inst_req_1;
      type_cast_1646_inst_ack_1<= rack(0);
      type_cast_1646_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1646_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc104x_xinput_dim0x_x2_1604,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1646_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1527_index_1_rename
    process(R_idxprom_1526_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1526_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1526_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1527_index_1_resize
    process(idxprom_1522) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1522;
      ov := iv(13 downto 0);
      R_idxprom_1526_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1527_root_address_inst
    process(array_obj_ref_1527_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1527_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1527_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1548_index_1_rename
    process(R_idxprom80_1547_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom80_1547_resized;
      ov(13 downto 0) := iv;
      R_idxprom80_1547_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1548_index_1_resize
    process(idxprom80_1543) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom80_1543;
      ov := iv(13 downto 0);
      R_idxprom80_1547_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1548_root_address_inst
    process(array_obj_ref_1548_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1548_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1548_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1532_addr_0
    process(ptr_deref_1532_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1532_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1532_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1532_base_resize
    process(arrayidx76_1529) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx76_1529;
      ov := iv(13 downto 0);
      ptr_deref_1532_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1532_gather_scatter
    process(ptr_deref_1532_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1532_data_0;
      ov(63 downto 0) := iv;
      tmp77_1533 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1532_root_address_inst
    process(ptr_deref_1532_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1532_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1532_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1552_addr_0
    process(ptr_deref_1552_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1552_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1552_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1552_base_resize
    process(arrayidx81_1550) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx81_1550;
      ov := iv(13 downto 0);
      ptr_deref_1552_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1552_gather_scatter
    process(tmp77_1533) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp77_1533;
      ov(63 downto 0) := iv;
      ptr_deref_1552_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1552_root_address_inst
    process(ptr_deref_1552_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1552_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1552_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1566_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1565;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1566_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1566_branch_req_0,
          ack0 => if_stmt_1566_branch_ack_0,
          ack1 => if_stmt_1566_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1621_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp111_1620;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1621_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1621_branch_req_0,
          ack0 => if_stmt_1621_branch_ack_0,
          ack1 => if_stmt_1621_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1577_inst
    process(input_dim2x_x1_1415) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1415, type_cast_1576_wire_constant, tmp_var);
      add92_1578 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1585_inst
    process(input_dim1x_x1_1423) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1423, type_cast_1584_wire_constant, tmp_var);
      inc_1586 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1603_inst
    process(inc104_1599, input_dim0x_x2_1430) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc104_1599, input_dim0x_x2_1430, tmp_var);
      inc104x_xinput_dim0x_x2_1604 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1352_inst
    process(call10_1316) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call10_1316, type_cast_1351_wire_constant, tmp_var);
      add_1353 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1363_inst
    process(call13_1319) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call13_1319, type_cast_1362_wire_constant, tmp_var);
      add53_1364 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1447_inst
    process(call23_1331, tmp1_1443) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call23_1331, tmp1_1443, tmp_var);
      add_src_0x_x0_1448 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1461_inst
    process(sub_1358, mul_1457) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1358, mul_1457, tmp_var);
      sub43_1462 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1475_inst
    process(sub56_1369, mul49_1471) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub56_1369, mul49_1471, tmp_var);
      sub57_1476 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1501_inst
    process(mul71_1497, conv65_1486) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul71_1497, conv65_1486, tmp_var);
      add72_1502 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1511_inst
    process(mul73_1507, conv60_1480) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul73_1507, conv60_1480, tmp_var);
      add74_1512 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1559_inst
    process(conv60_1480) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv60_1480, type_cast_1558_wire_constant, tmp_var);
      add85_1560 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1652_inst
    process(indvar_1408) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1408, type_cast_1651_wire_constant, tmp_var);
      indvarx_xnext_1653 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1346_inst
    process(call19_1325) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call19_1325, type_cast_1345_wire_constant, tmp_var);
      conv37_1347 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1374_inst
    process(call30_1340) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call30_1340, type_cast_1373_wire_constant, tmp_var);
      conv63_1375 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1380_inst
    process(call27_1337) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call27_1337, type_cast_1379_wire_constant, tmp_var);
      conv68_1381 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1386_inst
    process(call4_1310) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call4_1310, type_cast_1385_wire_constant, tmp_var);
      conv88_1387 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1392_inst
    process(call1_1307) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call1_1307, type_cast_1391_wire_constant, tmp_var);
      conv99_1393 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1404_inst
    process(conv109_1399) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv109_1399, type_cast_1403_wire_constant, tmp_var);
      shr110125_1405 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1485_inst
    process(sub57_1476) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(sub57_1476, type_cast_1484_wire_constant, tmp_var);
      conv65_1486 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1491_inst
    process(sub43_1462) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(sub43_1462, type_cast_1490_wire_constant, tmp_var);
      conv70_1492 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1594_inst
    process(conv96_1590, conv99_1393) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv96_1590, conv99_1393, tmp_var);
      cmp100_1595 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1619_inst
    process(conv106_1615, shr110125_1405) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv106_1615, shr110125_1405, tmp_var);
      cmp111_1620 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1398_inst
    process(call_1304) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1304, type_cast_1397_wire_constant, tmp_var);
      conv109_1399 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1517_inst
    process(add_src_0x_x0_1448) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_1448, type_cast_1516_wire_constant, tmp_var);
      shr_1518 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1538_inst
    process(add74_1512) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add74_1512, type_cast_1537_wire_constant, tmp_var);
      shr79_1539 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1442_inst
    process(indvar_1408) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1408, type_cast_1441_wire_constant, tmp_var);
      tmp1_1443 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1456_inst
    process(conv35_1452, conv37_1347) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv35_1452, conv37_1347, tmp_var);
      mul_1457 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1470_inst
    process(conv46_1466, conv37_1347) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv46_1466, conv37_1347, tmp_var);
      mul49_1471 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1496_inst
    process(conv70_1492, conv68_1381) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv70_1492, conv68_1381, tmp_var);
      mul71_1497 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1506_inst
    process(add72_1502, conv63_1375) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add72_1502, conv63_1375, tmp_var);
      mul73_1507 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1357_inst
    process(add_1353, call21_1328) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add_1353, call21_1328, tmp_var);
      sub_1358 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1368_inst
    process(add53_1364, call21_1328) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add53_1364, call21_1328, tmp_var);
      sub56_1369 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1564_inst
    process(add85_1560, conv88_1387) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add85_1560, conv88_1387, tmp_var);
      cmp_1565 <= tmp_var; --
    end process;
    -- shared split operator group (33) : array_obj_ref_1527_index_offset 
    ApIntAdd_group_33: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1526_scaled;
      array_obj_ref_1527_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1527_index_offset_req_0;
      array_obj_ref_1527_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1527_index_offset_req_1;
      array_obj_ref_1527_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_33_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_33_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_33",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : array_obj_ref_1548_index_offset 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom80_1547_scaled;
      array_obj_ref_1548_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1548_index_offset_req_0;
      array_obj_ref_1548_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1548_index_offset_req_1;
      array_obj_ref_1548_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared load operator group (0) : ptr_deref_1532_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1532_load_0_req_0;
      ptr_deref_1532_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1532_load_0_req_1;
      ptr_deref_1532_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1532_word_address_0;
      ptr_deref_1532_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1552_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1552_store_0_req_0;
      ptr_deref_1552_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1552_store_0_req_1;
      ptr_deref_1552_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1552_word_address_0;
      data_in <= ptr_deref_1552_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1339_inst RPIPE_Block0_start_1336_inst RPIPE_Block0_start_1333_inst RPIPE_Block0_start_1330_inst RPIPE_Block0_start_1327_inst RPIPE_Block0_start_1324_inst RPIPE_Block0_start_1321_inst RPIPE_Block0_start_1318_inst RPIPE_Block0_start_1315_inst RPIPE_Block0_start_1312_inst RPIPE_Block0_start_1309_inst RPIPE_Block0_start_1306_inst RPIPE_Block0_start_1303_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(415 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 12 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 12 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 12 downto 0);
      signal guard_vector : std_logic_vector( 12 downto 0);
      constant outBUFs : IntegerArray(12 downto 0) := (12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(12 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false);
      constant guardBuffering: IntegerArray(12 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2);
      -- 
    begin -- 
      reqL_unguarded(12) <= RPIPE_Block0_start_1339_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block0_start_1336_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block0_start_1333_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block0_start_1330_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block0_start_1327_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block0_start_1324_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block0_start_1321_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_start_1318_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_start_1315_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_start_1312_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_start_1309_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_start_1306_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_start_1303_inst_req_0;
      RPIPE_Block0_start_1339_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block0_start_1336_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block0_start_1333_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block0_start_1330_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block0_start_1327_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block0_start_1324_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block0_start_1321_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_start_1318_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_start_1315_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_start_1312_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_start_1309_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_start_1306_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_start_1303_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(12) <= RPIPE_Block0_start_1339_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block0_start_1336_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block0_start_1333_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block0_start_1330_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block0_start_1327_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block0_start_1324_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block0_start_1321_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_start_1318_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_start_1315_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_start_1312_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_start_1309_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_start_1306_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_start_1303_inst_req_1;
      RPIPE_Block0_start_1339_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block0_start_1336_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block0_start_1333_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block0_start_1330_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block0_start_1327_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block0_start_1324_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block0_start_1321_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_start_1318_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_start_1315_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_start_1312_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_start_1309_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_start_1306_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_start_1303_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      call30_1340 <= data_out(415 downto 384);
      call27_1337 <= data_out(383 downto 352);
      call24_1334 <= data_out(351 downto 320);
      call23_1331 <= data_out(319 downto 288);
      call21_1328 <= data_out(287 downto 256);
      call19_1325 <= data_out(255 downto 224);
      call16_1322 <= data_out(223 downto 192);
      call13_1319 <= data_out(191 downto 160);
      call10_1316 <= data_out(159 downto 128);
      call7_1313 <= data_out(127 downto 96);
      call4_1310 <= data_out(95 downto 64);
      call1_1307 <= data_out(63 downto 32);
      call_1304 <= data_out(31 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 13, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 32,  num_reqs => 13,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1657_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1657_inst_req_0;
      WPIPE_Block0_done_1657_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1657_inst_req_1;
      WPIPE_Block0_done_1657_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1659_wire_constant;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(31 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_4179_start: Boolean;
  signal convTransposeB_CP_4179_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_Block1_start_1677_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1689_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1674_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1671_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1683_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1686_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1674_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1677_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1689_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1683_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1692_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1701_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1683_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1683_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1692_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1692_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1686_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1701_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1677_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1695_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1668_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1701_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1677_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1668_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1695_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1692_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1686_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1695_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1668_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1686_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1680_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1695_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1668_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1671_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1674_inst_req_1 : boolean;
  signal type_cast_1721_inst_req_0 : boolean;
  signal type_cast_1721_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1674_inst_ack_1 : boolean;
  signal type_cast_1900_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1704_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1698_inst_ack_1 : boolean;
  signal type_cast_1900_inst_req_0 : boolean;
  signal type_cast_1900_inst_ack_0 : boolean;
  signal type_cast_1900_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1704_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1698_inst_req_1 : boolean;
  signal type_cast_1858_inst_req_1 : boolean;
  signal type_cast_1858_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1704_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1698_inst_ack_0 : boolean;
  signal type_cast_1858_inst_req_0 : boolean;
  signal type_cast_1858_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1704_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1698_inst_req_0 : boolean;
  signal array_obj_ref_1906_index_offset_req_0 : boolean;
  signal array_obj_ref_1906_index_offset_ack_0 : boolean;
  signal type_cast_1830_inst_req_1 : boolean;
  signal type_cast_1830_inst_ack_1 : boolean;
  signal type_cast_1721_inst_req_1 : boolean;
  signal type_cast_1721_inst_ack_1 : boolean;
  signal array_obj_ref_1906_index_offset_req_1 : boolean;
  signal array_obj_ref_1906_index_offset_ack_1 : boolean;
  signal type_cast_1830_inst_req_0 : boolean;
  signal type_cast_1830_inst_ack_0 : boolean;
  signal addr_of_1907_final_reg_req_0 : boolean;
  signal addr_of_1907_final_reg_ack_0 : boolean;
  signal RPIPE_Block1_start_1701_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1680_inst_req_1 : boolean;
  signal type_cast_1844_inst_req_0 : boolean;
  signal type_cast_1844_inst_ack_0 : boolean;
  signal type_cast_1844_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1689_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1671_inst_ack_1 : boolean;
  signal RPIPE_Block1_start_1689_inst_req_0 : boolean;
  signal type_cast_1844_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1671_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1680_inst_ack_0 : boolean;
  signal addr_of_1907_final_reg_req_1 : boolean;
  signal addr_of_1907_final_reg_ack_1 : boolean;
  signal RPIPE_Block1_start_1680_inst_req_0 : boolean;
  signal ptr_deref_1911_load_0_req_0 : boolean;
  signal ptr_deref_1911_load_0_ack_0 : boolean;
  signal ptr_deref_1911_load_0_req_1 : boolean;
  signal ptr_deref_1911_load_0_ack_1 : boolean;
  signal type_cast_1921_inst_req_0 : boolean;
  signal type_cast_1921_inst_ack_0 : boolean;
  signal type_cast_1921_inst_req_1 : boolean;
  signal type_cast_1921_inst_ack_1 : boolean;
  signal array_obj_ref_1927_index_offset_req_0 : boolean;
  signal array_obj_ref_1927_index_offset_ack_0 : boolean;
  signal array_obj_ref_1927_index_offset_req_1 : boolean;
  signal array_obj_ref_1927_index_offset_ack_1 : boolean;
  signal addr_of_1928_final_reg_req_0 : boolean;
  signal addr_of_1928_final_reg_ack_0 : boolean;
  signal addr_of_1928_final_reg_req_1 : boolean;
  signal addr_of_1928_final_reg_ack_1 : boolean;
  signal ptr_deref_1931_store_0_req_0 : boolean;
  signal ptr_deref_1931_store_0_ack_0 : boolean;
  signal ptr_deref_1931_store_0_req_1 : boolean;
  signal ptr_deref_1931_store_0_ack_1 : boolean;
  signal if_stmt_1945_branch_req_0 : boolean;
  signal if_stmt_1945_branch_ack_1 : boolean;
  signal if_stmt_1945_branch_ack_0 : boolean;
  signal type_cast_1968_inst_req_0 : boolean;
  signal type_cast_1968_inst_ack_0 : boolean;
  signal type_cast_1968_inst_req_1 : boolean;
  signal type_cast_1968_inst_ack_1 : boolean;
  signal type_cast_1977_inst_req_0 : boolean;
  signal type_cast_1977_inst_ack_0 : boolean;
  signal type_cast_1977_inst_req_1 : boolean;
  signal type_cast_1977_inst_ack_1 : boolean;
  signal type_cast_1993_inst_req_0 : boolean;
  signal type_cast_1993_inst_ack_0 : boolean;
  signal type_cast_1993_inst_req_1 : boolean;
  signal type_cast_1993_inst_ack_1 : boolean;
  signal if_stmt_2000_branch_req_0 : boolean;
  signal if_stmt_2000_branch_ack_1 : boolean;
  signal if_stmt_2000_branch_ack_0 : boolean;
  signal WPIPE_Block1_done_2036_inst_req_0 : boolean;
  signal WPIPE_Block1_done_2036_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2036_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2036_inst_ack_1 : boolean;
  signal type_cast_1815_inst_req_0 : boolean;
  signal type_cast_1815_inst_ack_0 : boolean;
  signal type_cast_1815_inst_req_1 : boolean;
  signal type_cast_1815_inst_ack_1 : boolean;
  signal phi_stmt_1810_req_1 : boolean;
  signal phi_stmt_1803_req_0 : boolean;
  signal phi_stmt_1796_req_1 : boolean;
  signal phi_stmt_1789_req_1 : boolean;
  signal type_cast_1813_inst_req_0 : boolean;
  signal type_cast_1813_inst_ack_0 : boolean;
  signal type_cast_1813_inst_req_1 : boolean;
  signal type_cast_1813_inst_ack_1 : boolean;
  signal phi_stmt_1810_req_0 : boolean;
  signal type_cast_1809_inst_req_0 : boolean;
  signal type_cast_1809_inst_ack_0 : boolean;
  signal type_cast_1809_inst_req_1 : boolean;
  signal type_cast_1809_inst_ack_1 : boolean;
  signal phi_stmt_1803_req_1 : boolean;
  signal type_cast_1799_inst_req_0 : boolean;
  signal type_cast_1799_inst_ack_0 : boolean;
  signal type_cast_1799_inst_req_1 : boolean;
  signal type_cast_1799_inst_ack_1 : boolean;
  signal phi_stmt_1796_req_0 : boolean;
  signal type_cast_1792_inst_req_0 : boolean;
  signal type_cast_1792_inst_ack_0 : boolean;
  signal type_cast_1792_inst_req_1 : boolean;
  signal type_cast_1792_inst_ack_1 : boolean;
  signal phi_stmt_1789_req_0 : boolean;
  signal phi_stmt_1789_ack_0 : boolean;
  signal phi_stmt_1796_ack_0 : boolean;
  signal phi_stmt_1803_ack_0 : boolean;
  signal phi_stmt_1810_ack_0 : boolean;
  signal type_cast_2023_inst_req_0 : boolean;
  signal type_cast_2023_inst_ack_0 : boolean;
  signal type_cast_2023_inst_req_1 : boolean;
  signal type_cast_2023_inst_ack_1 : boolean;
  signal phi_stmt_2020_req_0 : boolean;
  signal type_cast_2017_inst_req_0 : boolean;
  signal type_cast_2017_inst_ack_0 : boolean;
  signal type_cast_2017_inst_req_1 : boolean;
  signal type_cast_2017_inst_ack_1 : boolean;
  signal phi_stmt_2014_req_0 : boolean;
  signal phi_stmt_2007_req_0 : boolean;
  signal type_cast_2025_inst_req_0 : boolean;
  signal type_cast_2025_inst_ack_0 : boolean;
  signal type_cast_2025_inst_req_1 : boolean;
  signal type_cast_2025_inst_ack_1 : boolean;
  signal phi_stmt_2020_req_1 : boolean;
  signal type_cast_2019_inst_req_0 : boolean;
  signal type_cast_2019_inst_ack_0 : boolean;
  signal type_cast_2019_inst_req_1 : boolean;
  signal type_cast_2019_inst_ack_1 : boolean;
  signal phi_stmt_2014_req_1 : boolean;
  signal type_cast_2013_inst_req_0 : boolean;
  signal type_cast_2013_inst_ack_0 : boolean;
  signal type_cast_2013_inst_req_1 : boolean;
  signal type_cast_2013_inst_ack_1 : boolean;
  signal phi_stmt_2007_req_1 : boolean;
  signal phi_stmt_2007_ack_0 : boolean;
  signal phi_stmt_2014_ack_0 : boolean;
  signal phi_stmt_2020_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_4179_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4179_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_4179_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_4179_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_4179: Block -- control-path 
    signal convTransposeB_CP_4179_elements: BooleanArray(115 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_4179_elements(0) <= convTransposeB_CP_4179_start;
    convTransposeB_CP_4179_symbol <= convTransposeB_CP_4179_elements(66);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705__entry__
      -- CP-element group 0: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1668_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/$entry
      -- CP-element group 0: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1668_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1666/branch_block_stmt_1666__entry__
      -- CP-element group 0: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1668_Sample/rr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1666/$entry
      -- 
    rr_4227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(0), ack => RPIPE_Block1_start_1668_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	115 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	77 
    -- CP-element group 1: 	74 
    -- CP-element group 1: 	75 
    -- CP-element group 1: 	78 
    -- CP-element group 1: 	80 
    -- CP-element group 1: 	81 
    -- CP-element group 1: 	83 
    -- CP-element group 1: 	84 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_1666/assign_stmt_2032__exit__
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_1666/merge_stmt_2006__exit__
      -- CP-element group 1: 	 branch_block_stmt_1666/assign_stmt_2032__entry__
      -- CP-element group 1: 	 branch_block_stmt_1666/assign_stmt_2032/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/assign_stmt_2032/$exit
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1810/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1813/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1813/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1813/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1813/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1813/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1813/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1803/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1796/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1789/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_sources/type_cast_1792/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_sources/type_cast_1792/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_sources/type_cast_1792/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_sources/type_cast_1792/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_sources/type_cast_1792/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_sources/type_cast_1792/SplitProtocol/Update/cr
      -- 
    rr_4858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(1), ack => type_cast_1813_inst_req_0); -- 
    cr_4863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(1), ack => type_cast_1813_inst_req_1); -- 
    rr_4881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(1), ack => type_cast_1809_inst_req_0); -- 
    cr_4886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(1), ack => type_cast_1809_inst_req_1); -- 
    rr_4904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(1), ack => type_cast_1799_inst_req_0); -- 
    cr_4909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(1), ack => type_cast_1799_inst_req_1); -- 
    rr_4927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(1), ack => type_cast_1792_inst_req_0); -- 
    cr_4932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(1), ack => type_cast_1792_inst_req_1); -- 
    convTransposeB_CP_4179_elements(1) <= convTransposeB_CP_4179_elements(115);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1668_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1668_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1668_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1668_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1668_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1668_Update/cr
      -- 
    ra_4228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1668_inst_ack_0, ack => convTransposeB_CP_4179_elements(2)); -- 
    cr_4232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(2), ack => RPIPE_Block1_start_1668_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1668_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1668_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1668_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1671_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1671_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1671_Sample/rr
      -- 
    ca_4233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1668_inst_ack_1, ack => convTransposeB_CP_4179_elements(3)); -- 
    rr_4241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(3), ack => RPIPE_Block1_start_1671_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1671_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1671_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1671_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1671_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1671_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1671_Update/$entry
      -- 
    ra_4242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1671_inst_ack_0, ack => convTransposeB_CP_4179_elements(4)); -- 
    cr_4246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(4), ack => RPIPE_Block1_start_1671_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1671_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1674_Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1674_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1674_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1671_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1671_Update/$exit
      -- 
    ca_4247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1671_inst_ack_1, ack => convTransposeB_CP_4179_elements(5)); -- 
    rr_4255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(5), ack => RPIPE_Block1_start_1674_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1674_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1674_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1674_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1674_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1674_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1674_sample_completed_
      -- 
    ra_4256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1674_inst_ack_0, ack => convTransposeB_CP_4179_elements(6)); -- 
    cr_4260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(6), ack => RPIPE_Block1_start_1674_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1677_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1677_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1677_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1674_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1674_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1674_update_completed_
      -- 
    ca_4261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1674_inst_ack_1, ack => convTransposeB_CP_4179_elements(7)); -- 
    rr_4269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(7), ack => RPIPE_Block1_start_1677_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1677_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1677_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1677_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1677_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1677_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1677_Update/cr
      -- 
    ra_4270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1677_inst_ack_0, ack => convTransposeB_CP_4179_elements(8)); -- 
    cr_4274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(8), ack => RPIPE_Block1_start_1677_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1677_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1677_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1677_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1680_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1680_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1680_Sample/rr
      -- 
    ca_4275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1677_inst_ack_1, ack => convTransposeB_CP_4179_elements(9)); -- 
    rr_4283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(9), ack => RPIPE_Block1_start_1680_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1680_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1680_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1680_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1680_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1680_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1680_Sample/ra
      -- 
    ra_4284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1680_inst_ack_0, ack => convTransposeB_CP_4179_elements(10)); -- 
    cr_4288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(10), ack => RPIPE_Block1_start_1680_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1683_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1683_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1683_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1680_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1680_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1680_Update/$exit
      -- 
    ca_4289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1680_inst_ack_1, ack => convTransposeB_CP_4179_elements(11)); -- 
    rr_4297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(11), ack => RPIPE_Block1_start_1683_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1683_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1683_Update/cr
      -- CP-element group 12: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1683_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1683_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1683_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1683_Sample/$exit
      -- 
    ra_4298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1683_inst_ack_0, ack => convTransposeB_CP_4179_elements(12)); -- 
    cr_4302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(12), ack => RPIPE_Block1_start_1683_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1686_Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1683_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1686_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1683_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1683_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1686_sample_start_
      -- 
    ca_4303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1683_inst_ack_1, ack => convTransposeB_CP_4179_elements(13)); -- 
    rr_4311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(13), ack => RPIPE_Block1_start_1686_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1686_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1686_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1686_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1686_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1686_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1686_update_start_
      -- 
    ra_4312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1686_inst_ack_0, ack => convTransposeB_CP_4179_elements(14)); -- 
    cr_4316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(14), ack => RPIPE_Block1_start_1686_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1686_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1686_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1686_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1689_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1689_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1689_Sample/$entry
      -- 
    ca_4317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1686_inst_ack_1, ack => convTransposeB_CP_4179_elements(15)); -- 
    rr_4325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(15), ack => RPIPE_Block1_start_1689_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1689_Update/cr
      -- CP-element group 16: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1689_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1689_update_start_
      -- CP-element group 16: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1689_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1689_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1689_Sample/$exit
      -- 
    ra_4326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1689_inst_ack_0, ack => convTransposeB_CP_4179_elements(16)); -- 
    cr_4330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(16), ack => RPIPE_Block1_start_1689_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1692_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1689_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1689_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1692_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1689_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1692_Sample/$entry
      -- 
    ca_4331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1689_inst_ack_1, ack => convTransposeB_CP_4179_elements(17)); -- 
    rr_4339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(17), ack => RPIPE_Block1_start_1692_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1692_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1692_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1692_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1692_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1692_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1692_Sample/$exit
      -- 
    ra_4340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1692_inst_ack_0, ack => convTransposeB_CP_4179_elements(18)); -- 
    cr_4344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(18), ack => RPIPE_Block1_start_1692_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1692_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1692_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1692_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1695_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1695_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1695_Sample/rr
      -- 
    ca_4345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1692_inst_ack_1, ack => convTransposeB_CP_4179_elements(19)); -- 
    rr_4353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(19), ack => RPIPE_Block1_start_1695_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1695_update_start_
      -- CP-element group 20: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1695_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1695_Update/cr
      -- CP-element group 20: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1695_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1695_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1695_Sample/ra
      -- 
    ra_4354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1695_inst_ack_0, ack => convTransposeB_CP_4179_elements(20)); -- 
    cr_4358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(20), ack => RPIPE_Block1_start_1695_inst_req_1); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1695_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1695_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1695_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1698_Sample/rr
      -- CP-element group 21: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1698_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1698_sample_start_
      -- 
    ca_4359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1695_inst_ack_1, ack => convTransposeB_CP_4179_elements(21)); -- 
    rr_4367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(21), ack => RPIPE_Block1_start_1698_inst_req_0); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1698_Update/cr
      -- CP-element group 22: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1698_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1698_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1698_update_start_
      -- CP-element group 22: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1698_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1698_Update/$entry
      -- 
    ra_4368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1698_inst_ack_0, ack => convTransposeB_CP_4179_elements(22)); -- 
    cr_4372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(22), ack => RPIPE_Block1_start_1698_inst_req_1); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1698_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1701_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1701_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1701_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1698_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1698_Update/$exit
      -- 
    ca_4373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1698_inst_ack_1, ack => convTransposeB_CP_4179_elements(23)); -- 
    rr_4381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(23), ack => RPIPE_Block1_start_1701_inst_req_0); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1701_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1701_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1701_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1701_Update/cr
      -- CP-element group 24: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1701_update_start_
      -- CP-element group 24: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1701_sample_completed_
      -- 
    ra_4382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1701_inst_ack_0, ack => convTransposeB_CP_4179_elements(24)); -- 
    cr_4386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(24), ack => RPIPE_Block1_start_1701_inst_req_1); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1701_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1701_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1704_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1704_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1704_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1701_Update/ca
      -- 
    ca_4387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1701_inst_ack_1, ack => convTransposeB_CP_4179_elements(25)); -- 
    rr_4395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(25), ack => RPIPE_Block1_start_1704_inst_req_0); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1704_Update/cr
      -- CP-element group 26: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1704_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1704_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1704_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1704_update_start_
      -- CP-element group 26: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1704_sample_completed_
      -- 
    ra_4396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1704_inst_ack_0, ack => convTransposeB_CP_4179_elements(26)); -- 
    cr_4400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(26), ack => RPIPE_Block1_start_1704_inst_req_1); -- 
    -- CP-element group 27:  fork  transition  place  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (13) 
      -- CP-element group 27: 	 branch_block_stmt_1666/assign_stmt_1712_to_assign_stmt_1786__entry__
      -- CP-element group 27: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705__exit__
      -- CP-element group 27: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1704_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1666/assign_stmt_1712_to_assign_stmt_1786/type_cast_1721_update_start_
      -- CP-element group 27: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/$exit
      -- CP-element group 27: 	 branch_block_stmt_1666/assign_stmt_1712_to_assign_stmt_1786/type_cast_1721_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_1666/assign_stmt_1712_to_assign_stmt_1786/type_cast_1721_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1666/assign_stmt_1712_to_assign_stmt_1786/type_cast_1721_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1666/assign_stmt_1712_to_assign_stmt_1786/$entry
      -- CP-element group 27: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1704_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1666/assign_stmt_1669_to_assign_stmt_1705/RPIPE_Block1_start_1704_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1666/assign_stmt_1712_to_assign_stmt_1786/type_cast_1721_Update/cr
      -- CP-element group 27: 	 branch_block_stmt_1666/assign_stmt_1712_to_assign_stmt_1786/type_cast_1721_Update/$entry
      -- 
    ca_4401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1704_inst_ack_1, ack => convTransposeB_CP_4179_elements(27)); -- 
    rr_4412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(27), ack => type_cast_1721_inst_req_0); -- 
    cr_4417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(27), ack => type_cast_1721_inst_req_1); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1666/assign_stmt_1712_to_assign_stmt_1786/type_cast_1721_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1666/assign_stmt_1712_to_assign_stmt_1786/type_cast_1721_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1666/assign_stmt_1712_to_assign_stmt_1786/type_cast_1721_Sample/ra
      -- 
    ra_4413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1721_inst_ack_0, ack => convTransposeB_CP_4179_elements(28)); -- 
    -- CP-element group 29:  fork  transition  place  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	67 
    -- CP-element group 29: 	68 
    -- CP-element group 29: 	72 
    -- CP-element group 29: 	70 
    -- CP-element group 29: 	71 
    -- CP-element group 29:  members (21) 
      -- CP-element group 29: 	 branch_block_stmt_1666/assign_stmt_1712_to_assign_stmt_1786__exit__
      -- CP-element group 29: 	 branch_block_stmt_1666/entry_whilex_xbody
      -- CP-element group 29: 	 branch_block_stmt_1666/assign_stmt_1712_to_assign_stmt_1786/type_cast_1721_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1666/assign_stmt_1712_to_assign_stmt_1786/$exit
      -- CP-element group 29: 	 branch_block_stmt_1666/assign_stmt_1712_to_assign_stmt_1786/type_cast_1721_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1666/assign_stmt_1712_to_assign_stmt_1786/type_cast_1721_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 29: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1810/$entry
      -- CP-element group 29: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1815/$entry
      -- CP-element group 29: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1815/SplitProtocol/$entry
      -- CP-element group 29: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1815/SplitProtocol/Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1815/SplitProtocol/Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1815/SplitProtocol/Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1815/SplitProtocol/Update/cr
      -- CP-element group 29: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1803/$entry
      -- CP-element group 29: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1796/$entry
      -- CP-element group 29: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1789/$entry
      -- CP-element group 29: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_sources/$entry
      -- 
    ca_4418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1721_inst_ack_1, ack => convTransposeB_CP_4179_elements(29)); -- 
    rr_4808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(29), ack => type_cast_1815_inst_req_0); -- 
    cr_4813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(29), ack => type_cast_1815_inst_req_1); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	92 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1830_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1830_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1830_Sample/ra
      -- 
    ra_4430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1830_inst_ack_0, ack => convTransposeB_CP_4179_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	92 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	44 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1830_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1830_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1830_Update/$exit
      -- 
    ca_4435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1830_inst_ack_1, ack => convTransposeB_CP_4179_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	92 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1844_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1844_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1844_Sample/$exit
      -- 
    ra_4444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1844_inst_ack_0, ack => convTransposeB_CP_4179_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	92 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	44 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1844_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1844_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1844_Update/$exit
      -- 
    ca_4449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1844_inst_ack_1, ack => convTransposeB_CP_4179_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	92 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1858_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1858_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1858_Sample/$exit
      -- 
    ra_4458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1858_inst_ack_0, ack => convTransposeB_CP_4179_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	92 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	44 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1858_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1858_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1858_update_completed_
      -- 
    ca_4463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1858_inst_ack_1, ack => convTransposeB_CP_4179_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	92 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1900_Sample/ra
      -- CP-element group 36: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1900_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1900_sample_completed_
      -- 
    ra_4472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1900_inst_ack_0, ack => convTransposeB_CP_4179_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	92 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (16) 
      -- CP-element group 37: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_index_scale_1/$entry
      -- CP-element group 37: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_index_scale_1/$exit
      -- CP-element group 37: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_index_scale_1/scale_rename_req
      -- CP-element group 37: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_index_resized_1
      -- CP-element group 37: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_index_scaled_1
      -- CP-element group 37: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_index_computed_1
      -- CP-element group 37: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_index_scale_1/scale_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1900_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1900_Update/ca
      -- CP-element group 37: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1900_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_index_resize_1/index_resize_req
      -- CP-element group 37: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_index_resize_1/index_resize_ack
      -- CP-element group 37: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_index_resize_1/$entry
      -- CP-element group 37: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_index_resize_1/$exit
      -- CP-element group 37: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_final_index_sum_regn_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_final_index_sum_regn_Sample/req
      -- 
    ca_4477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1900_inst_ack_1, ack => convTransposeB_CP_4179_elements(37)); -- 
    req_4502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(37), ack => array_obj_ref_1906_index_offset_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	54 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_final_index_sum_regn_sample_complete
      -- CP-element group 38: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_final_index_sum_regn_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_final_index_sum_regn_Sample/ack
      -- 
    ack_4503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1906_index_offset_ack_0, ack => convTransposeB_CP_4179_elements(38)); -- 
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	92 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (11) 
      -- CP-element group 39: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_offset_calculated
      -- CP-element group 39: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1907_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_final_index_sum_regn_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_final_index_sum_regn_Update/ack
      -- CP-element group 39: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1907_request/$entry
      -- CP-element group 39: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1907_request/req
      -- 
    ack_4508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1906_index_offset_ack_1, ack => convTransposeB_CP_4179_elements(39)); -- 
    req_4517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(39), ack => addr_of_1907_final_reg_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1907_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1907_request/$exit
      -- CP-element group 40: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1907_request/ack
      -- 
    ack_4518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1907_final_reg_ack_0, ack => convTransposeB_CP_4179_elements(40)); -- 
    -- CP-element group 41:  join  fork  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	92 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (24) 
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1907_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_base_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_word_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1907_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1907_complete/ack
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_base_address_resized
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_base_addr_resize/$entry
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_base_addr_resize/$exit
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_base_addr_resize/base_resize_req
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_base_addr_resize/base_resize_ack
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_base_plus_offset/$entry
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_base_plus_offset/$exit
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_word_addrgen/$entry
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_word_addrgen/$exit
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_word_addrgen/root_register_req
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_word_addrgen/root_register_ack
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Sample/word_access_start/$entry
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Sample/word_access_start/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Sample/word_access_start/word_0/rr
      -- 
    ack_4523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1907_final_reg_ack_1, ack => convTransposeB_CP_4179_elements(41)); -- 
    rr_4556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(41), ack => ptr_deref_1911_load_0_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Sample/word_access_start/$exit
      -- CP-element group 42: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Sample/word_access_start/word_0/$exit
      -- CP-element group 42: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Sample/word_access_start/word_0/ra
      -- 
    ra_4557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1911_load_0_ack_0, ack => convTransposeB_CP_4179_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	92 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	51 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Update/word_access_complete/$exit
      -- CP-element group 43: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Update/word_access_complete/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Update/word_access_complete/word_0/ca
      -- CP-element group 43: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Update/ptr_deref_1911_Merge/$entry
      -- CP-element group 43: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Update/ptr_deref_1911_Merge/$exit
      -- CP-element group 43: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Update/ptr_deref_1911_Merge/merge_req
      -- CP-element group 43: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Update/ptr_deref_1911_Merge/merge_ack
      -- 
    ca_4568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1911_load_0_ack_1, ack => convTransposeB_CP_4179_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	31 
    -- CP-element group 44: 	35 
    -- CP-element group 44: 	33 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1921_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1921_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1921_Sample/rr
      -- 
    rr_4581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(44), ack => type_cast_1921_inst_req_0); -- 
    convTransposeB_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(31) & convTransposeB_CP_4179_elements(35) & convTransposeB_CP_4179_elements(33);
      gj_convTransposeB_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1921_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1921_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1921_Sample/ra
      -- 
    ra_4582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1921_inst_ack_0, ack => convTransposeB_CP_4179_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	92 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (16) 
      -- CP-element group 46: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1921_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1921_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1921_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_index_resized_1
      -- CP-element group 46: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_index_scaled_1
      -- CP-element group 46: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_index_computed_1
      -- CP-element group 46: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_index_resize_1/$entry
      -- CP-element group 46: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_index_resize_1/$exit
      -- CP-element group 46: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_index_resize_1/index_resize_req
      -- CP-element group 46: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_index_resize_1/index_resize_ack
      -- CP-element group 46: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_index_scale_1/$entry
      -- CP-element group 46: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_index_scale_1/$exit
      -- CP-element group 46: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_index_scale_1/scale_rename_req
      -- CP-element group 46: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_index_scale_1/scale_rename_ack
      -- CP-element group 46: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_final_index_sum_regn_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_final_index_sum_regn_Sample/req
      -- 
    ca_4587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1921_inst_ack_1, ack => convTransposeB_CP_4179_elements(46)); -- 
    req_4612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(46), ack => array_obj_ref_1927_index_offset_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	54 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_final_index_sum_regn_sample_complete
      -- CP-element group 47: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_final_index_sum_regn_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_final_index_sum_regn_Sample/ack
      -- 
    ack_4613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1927_index_offset_ack_0, ack => convTransposeB_CP_4179_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	92 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (11) 
      -- CP-element group 48: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_root_address_calculated
      -- CP-element group 48: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1928_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_offset_calculated
      -- CP-element group 48: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_final_index_sum_regn_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_final_index_sum_regn_Update/ack
      -- CP-element group 48: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_base_plus_offset/$entry
      -- CP-element group 48: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_base_plus_offset/$exit
      -- CP-element group 48: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_base_plus_offset/sum_rename_req
      -- CP-element group 48: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_base_plus_offset/sum_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1928_request/$entry
      -- CP-element group 48: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1928_request/req
      -- 
    ack_4618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1927_index_offset_ack_1, ack => convTransposeB_CP_4179_elements(48)); -- 
    req_4627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(48), ack => addr_of_1928_final_reg_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1928_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1928_request/$exit
      -- CP-element group 49: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1928_request/ack
      -- 
    ack_4628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1928_final_reg_ack_0, ack => convTransposeB_CP_4179_elements(49)); -- 
    -- CP-element group 50:  fork  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	92 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (19) 
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1928_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1928_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1928_complete/ack
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_base_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_word_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_base_address_resized
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_base_addr_resize/$entry
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_base_addr_resize/$exit
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_base_addr_resize/base_resize_req
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_base_addr_resize/base_resize_ack
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_base_plus_offset/sum_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_word_addrgen/$entry
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_word_addrgen/$exit
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_word_addrgen/root_register_req
      -- CP-element group 50: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_word_addrgen/root_register_ack
      -- 
    ack_4633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1928_final_reg_ack_1, ack => convTransposeB_CP_4179_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: 	43 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Sample/ptr_deref_1931_Split/$entry
      -- CP-element group 51: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Sample/ptr_deref_1931_Split/$exit
      -- CP-element group 51: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Sample/ptr_deref_1931_Split/split_req
      -- CP-element group 51: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Sample/ptr_deref_1931_Split/split_ack
      -- CP-element group 51: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Sample/word_access_start/word_0/rr
      -- 
    rr_4671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(51), ack => ptr_deref_1931_store_0_req_0); -- 
    convTransposeB_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(50) & convTransposeB_CP_4179_elements(43);
      gj_convTransposeB_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Sample/word_access_start/word_0/ra
      -- 
    ra_4672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1931_store_0_ack_0, ack => convTransposeB_CP_4179_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	92 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Update/word_access_complete/word_0/ca
      -- 
    ca_4683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1931_store_0_ack_1, ack => convTransposeB_CP_4179_elements(53)); -- 
    -- CP-element group 54:  branch  join  transition  place  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	47 
    -- CP-element group 54: 	38 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (10) 
      -- CP-element group 54: 	 branch_block_stmt_1666/if_stmt_1945__entry__
      -- CP-element group 54: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944__exit__
      -- CP-element group 54: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/$exit
      -- CP-element group 54: 	 branch_block_stmt_1666/if_stmt_1945_dead_link/$entry
      -- CP-element group 54: 	 branch_block_stmt_1666/if_stmt_1945_eval_test/$entry
      -- CP-element group 54: 	 branch_block_stmt_1666/if_stmt_1945_eval_test/$exit
      -- CP-element group 54: 	 branch_block_stmt_1666/if_stmt_1945_eval_test/branch_req
      -- CP-element group 54: 	 branch_block_stmt_1666/R_cmp_1946_place
      -- CP-element group 54: 	 branch_block_stmt_1666/if_stmt_1945_if_link/$entry
      -- CP-element group 54: 	 branch_block_stmt_1666/if_stmt_1945_else_link/$entry
      -- 
    branch_req_4691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(54), ack => if_stmt_1945_branch_req_0); -- 
    convTransposeB_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(47) & convTransposeB_CP_4179_elements(38) & convTransposeB_CP_4179_elements(53);
      gj_convTransposeB_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	101 
    -- CP-element group 55: 	102 
    -- CP-element group 55: 	104 
    -- CP-element group 55: 	105 
    -- CP-element group 55: 	107 
    -- CP-element group 55: 	108 
    -- CP-element group 55:  members (40) 
      -- CP-element group 55: 	 branch_block_stmt_1666/assign_stmt_1957__entry__
      -- CP-element group 55: 	 branch_block_stmt_1666/merge_stmt_1951__exit__
      -- CP-element group 55: 	 branch_block_stmt_1666/assign_stmt_1957__exit__
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134
      -- CP-element group 55: 	 branch_block_stmt_1666/if_stmt_1945_if_link/$exit
      -- CP-element group 55: 	 branch_block_stmt_1666/if_stmt_1945_if_link/if_choice_transition
      -- CP-element group 55: 	 branch_block_stmt_1666/whilex_xbody_ifx_xthen
      -- CP-element group 55: 	 branch_block_stmt_1666/assign_stmt_1957/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/assign_stmt_1957/$exit
      -- CP-element group 55: 	 branch_block_stmt_1666/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 55: 	 branch_block_stmt_1666/merge_stmt_1951_PhiReqMerge
      -- CP-element group 55: 	 branch_block_stmt_1666/merge_stmt_1951_PhiAck/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/merge_stmt_1951_PhiAck/$exit
      -- CP-element group 55: 	 branch_block_stmt_1666/merge_stmt_1951_PhiAck/dummy
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2020/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2025/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2025/SplitProtocol/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2025/SplitProtocol/Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2025/SplitProtocol/Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2025/SplitProtocol/Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2025/SplitProtocol/Update/cr
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2014/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2019/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2019/SplitProtocol/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2019/SplitProtocol/Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2019/SplitProtocol/Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2019/SplitProtocol/Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2019/SplitProtocol/Update/cr
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2007/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_sources/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_sources/type_cast_2013/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_sources/type_cast_2013/SplitProtocol/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_sources/type_cast_2013/SplitProtocol/Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_sources/type_cast_2013/SplitProtocol/Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_sources/type_cast_2013/SplitProtocol/Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_sources/type_cast_2013/SplitProtocol/Update/cr
      -- 
    if_choice_transition_4696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1945_branch_ack_1, ack => convTransposeB_CP_4179_elements(55)); -- 
    rr_5042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(55), ack => type_cast_2025_inst_req_0); -- 
    cr_5047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(55), ack => type_cast_2025_inst_req_1); -- 
    rr_5065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(55), ack => type_cast_2019_inst_req_0); -- 
    cr_5070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(55), ack => type_cast_2019_inst_req_1); -- 
    rr_5088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(55), ack => type_cast_2013_inst_req_0); -- 
    cr_5093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(55), ack => type_cast_2013_inst_req_1); -- 
    -- CP-element group 56:  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	62 
    -- CP-element group 56: 	60 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (24) 
      -- CP-element group 56: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999__entry__
      -- CP-element group 56: 	 branch_block_stmt_1666/merge_stmt_1959__exit__
      -- CP-element group 56: 	 branch_block_stmt_1666/if_stmt_1945_else_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_1666/if_stmt_1945_else_link/else_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_1666/whilex_xbody_ifx_xelse
      -- CP-element group 56: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/$entry
      -- CP-element group 56: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1968_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1968_update_start_
      -- CP-element group 56: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1968_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1968_Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1968_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1968_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1977_update_start_
      -- CP-element group 56: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1977_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1977_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1993_update_start_
      -- CP-element group 56: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1993_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1993_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_1666/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1666/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_1666/merge_stmt_1959_PhiReqMerge
      -- CP-element group 56: 	 branch_block_stmt_1666/merge_stmt_1959_PhiAck/$entry
      -- CP-element group 56: 	 branch_block_stmt_1666/merge_stmt_1959_PhiAck/$exit
      -- CP-element group 56: 	 branch_block_stmt_1666/merge_stmt_1959_PhiAck/dummy
      -- 
    else_choice_transition_4700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1945_branch_ack_0, ack => convTransposeB_CP_4179_elements(56)); -- 
    rr_4716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(56), ack => type_cast_1968_inst_req_0); -- 
    cr_4721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(56), ack => type_cast_1968_inst_req_1); -- 
    cr_4735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(56), ack => type_cast_1977_inst_req_1); -- 
    cr_4749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(56), ack => type_cast_1993_inst_req_1); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1968_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1968_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1968_Sample/ra
      -- 
    ra_4717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1968_inst_ack_0, ack => convTransposeB_CP_4179_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1968_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1968_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1968_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1977_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1977_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1977_Sample/rr
      -- 
    ca_4722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1968_inst_ack_1, ack => convTransposeB_CP_4179_elements(58)); -- 
    rr_4730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(58), ack => type_cast_1977_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1977_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1977_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1977_Sample/ra
      -- 
    ra_4731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1977_inst_ack_0, ack => convTransposeB_CP_4179_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	56 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1977_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1977_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1977_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1993_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1993_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1993_Sample/rr
      -- 
    ca_4736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1977_inst_ack_1, ack => convTransposeB_CP_4179_elements(60)); -- 
    rr_4744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(60), ack => type_cast_1993_inst_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1993_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1993_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1993_Sample/ra
      -- 
    ra_4745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1993_inst_ack_0, ack => convTransposeB_CP_4179_elements(61)); -- 
    -- CP-element group 62:  branch  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	56 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (13) 
      -- CP-element group 62: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999__exit__
      -- CP-element group 62: 	 branch_block_stmt_1666/if_stmt_2000__entry__
      -- CP-element group 62: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/$exit
      -- CP-element group 62: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1993_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1993_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1666/assign_stmt_1965_to_assign_stmt_1999/type_cast_1993_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_1666/if_stmt_2000_dead_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_1666/if_stmt_2000_eval_test/$entry
      -- CP-element group 62: 	 branch_block_stmt_1666/if_stmt_2000_eval_test/$exit
      -- CP-element group 62: 	 branch_block_stmt_1666/if_stmt_2000_eval_test/branch_req
      -- CP-element group 62: 	 branch_block_stmt_1666/R_cmp123_2001_place
      -- CP-element group 62: 	 branch_block_stmt_1666/if_stmt_2000_if_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_1666/if_stmt_2000_else_link/$entry
      -- 
    ca_4750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1993_inst_ack_1, ack => convTransposeB_CP_4179_elements(62)); -- 
    branch_req_4758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(62), ack => if_stmt_2000_branch_req_0); -- 
    -- CP-element group 63:  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (15) 
      -- CP-element group 63: 	 branch_block_stmt_1666/merge_stmt_2034__exit__
      -- CP-element group 63: 	 branch_block_stmt_1666/assign_stmt_2039__entry__
      -- CP-element group 63: 	 branch_block_stmt_1666/if_stmt_2000_if_link/$exit
      -- CP-element group 63: 	 branch_block_stmt_1666/if_stmt_2000_if_link/if_choice_transition
      -- CP-element group 63: 	 branch_block_stmt_1666/ifx_xelse_whilex_xend
      -- CP-element group 63: 	 branch_block_stmt_1666/assign_stmt_2039/$entry
      -- CP-element group 63: 	 branch_block_stmt_1666/assign_stmt_2039/WPIPE_Block1_done_2036_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1666/assign_stmt_2039/WPIPE_Block1_done_2036_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1666/assign_stmt_2039/WPIPE_Block1_done_2036_Sample/req
      -- CP-element group 63: 	 branch_block_stmt_1666/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 63: 	 branch_block_stmt_1666/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 63: 	 branch_block_stmt_1666/merge_stmt_2034_PhiReqMerge
      -- CP-element group 63: 	 branch_block_stmt_1666/merge_stmt_2034_PhiAck/$entry
      -- CP-element group 63: 	 branch_block_stmt_1666/merge_stmt_2034_PhiAck/$exit
      -- CP-element group 63: 	 branch_block_stmt_1666/merge_stmt_2034_PhiAck/dummy
      -- 
    if_choice_transition_4763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2000_branch_ack_1, ack => convTransposeB_CP_4179_elements(63)); -- 
    req_4783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(63), ack => WPIPE_Block1_done_2036_inst_req_0); -- 
    -- CP-element group 64:  fork  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	93 
    -- CP-element group 64: 	94 
    -- CP-element group 64: 	96 
    -- CP-element group 64: 	97 
    -- CP-element group 64: 	99 
    -- CP-element group 64:  members (22) 
      -- CP-element group 64: 	 branch_block_stmt_1666/if_stmt_2000_else_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_1666/if_stmt_2000_else_link/else_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2020/$entry
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/$entry
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2023/$entry
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2023/SplitProtocol/$entry
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2023/SplitProtocol/Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2023/SplitProtocol/Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2023/SplitProtocol/Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2023/SplitProtocol/Update/cr
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2014/$entry
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/$entry
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/$entry
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/$entry
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/Update/cr
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2007/$entry
      -- CP-element group 64: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_sources/$entry
      -- 
    else_choice_transition_4767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2000_branch_ack_0, ack => convTransposeB_CP_4179_elements(64)); -- 
    rr_4985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(64), ack => type_cast_2023_inst_req_0); -- 
    cr_4990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(64), ack => type_cast_2023_inst_req_1); -- 
    rr_5008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(64), ack => type_cast_2017_inst_req_0); -- 
    cr_5013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(64), ack => type_cast_2017_inst_req_1); -- 
    -- CP-element group 65:  transition  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (6) 
      -- CP-element group 65: 	 branch_block_stmt_1666/assign_stmt_2039/WPIPE_Block1_done_2036_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_1666/assign_stmt_2039/WPIPE_Block1_done_2036_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1666/assign_stmt_2039/WPIPE_Block1_done_2036_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_1666/assign_stmt_2039/WPIPE_Block1_done_2036_Sample/ack
      -- CP-element group 65: 	 branch_block_stmt_1666/assign_stmt_2039/WPIPE_Block1_done_2036_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1666/assign_stmt_2039/WPIPE_Block1_done_2036_Update/req
      -- 
    ack_4784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2036_inst_ack_0, ack => convTransposeB_CP_4179_elements(65)); -- 
    req_4788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(65), ack => WPIPE_Block1_done_2036_inst_req_1); -- 
    -- CP-element group 66:  transition  place  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (16) 
      -- CP-element group 66: 	 branch_block_stmt_1666/merge_stmt_2041__exit__
      -- CP-element group 66: 	 branch_block_stmt_1666/$exit
      -- CP-element group 66: 	 branch_block_stmt_1666/return__
      -- CP-element group 66: 	 branch_block_stmt_1666/branch_block_stmt_1666__exit__
      -- CP-element group 66: 	 $exit
      -- CP-element group 66: 	 branch_block_stmt_1666/assign_stmt_2039__exit__
      -- CP-element group 66: 	 branch_block_stmt_1666/assign_stmt_2039/$exit
      -- CP-element group 66: 	 branch_block_stmt_1666/assign_stmt_2039/WPIPE_Block1_done_2036_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_1666/assign_stmt_2039/WPIPE_Block1_done_2036_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_1666/assign_stmt_2039/WPIPE_Block1_done_2036_Update/ack
      -- CP-element group 66: 	 branch_block_stmt_1666/return___PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_1666/return___PhiReq/$exit
      -- CP-element group 66: 	 branch_block_stmt_1666/merge_stmt_2041_PhiReqMerge
      -- CP-element group 66: 	 branch_block_stmt_1666/merge_stmt_2041_PhiAck/$entry
      -- CP-element group 66: 	 branch_block_stmt_1666/merge_stmt_2041_PhiAck/$exit
      -- CP-element group 66: 	 branch_block_stmt_1666/merge_stmt_2041_PhiAck/dummy
      -- 
    ack_4789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2036_inst_ack_1, ack => convTransposeB_CP_4179_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	29 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1815/SplitProtocol/Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1815/SplitProtocol/Sample/ra
      -- 
    ra_4809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1815_inst_ack_0, ack => convTransposeB_CP_4179_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	29 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1815/SplitProtocol/Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1815/SplitProtocol/Update/ca
      -- 
    ca_4814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1815_inst_ack_1, ack => convTransposeB_CP_4179_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	73 
    -- CP-element group 69:  members (5) 
      -- CP-element group 69: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1810/$exit
      -- CP-element group 69: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/$exit
      -- CP-element group 69: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1815/$exit
      -- CP-element group 69: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1815/SplitProtocol/$exit
      -- CP-element group 69: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_req
      -- 
    phi_stmt_1810_req_4815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1810_req_4815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(69), ack => phi_stmt_1810_req_1); -- 
    convTransposeB_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(67) & convTransposeB_CP_4179_elements(68);
      gj_convTransposeB_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  output  delay-element  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	29 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	73 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1803/$exit
      -- CP-element group 70: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/$exit
      -- CP-element group 70: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1807_konst_delay_trans
      -- CP-element group 70: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_req
      -- 
    phi_stmt_1803_req_4823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1803_req_4823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(70), ack => phi_stmt_1803_req_0); -- 
    -- Element group convTransposeB_CP_4179_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => convTransposeB_CP_4179_elements(29), ack => convTransposeB_CP_4179_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  transition  output  delay-element  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	29 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1796/$exit
      -- CP-element group 71: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/$exit
      -- CP-element group 71: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1802_konst_delay_trans
      -- CP-element group 71: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_req
      -- 
    phi_stmt_1796_req_4831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1796_req_4831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(71), ack => phi_stmt_1796_req_1); -- 
    -- Element group convTransposeB_CP_4179_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => convTransposeB_CP_4179_elements(29), ack => convTransposeB_CP_4179_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  transition  output  delay-element  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	29 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1789/$exit
      -- CP-element group 72: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_sources/$exit
      -- CP-element group 72: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_sources/type_cast_1795_konst_delay_trans
      -- CP-element group 72: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_req
      -- 
    phi_stmt_1789_req_4839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1789_req_4839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(72), ack => phi_stmt_1789_req_1); -- 
    -- Element group convTransposeB_CP_4179_elements(72) is a control-delay.
    cp_element_72_delay: control_delay_element  generic map(name => " 72_delay", delay_value => 1)  port map(req => convTransposeB_CP_4179_elements(29), ack => convTransposeB_CP_4179_elements(72), clk => clk, reset =>reset);
    -- CP-element group 73:  join  transition  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: 	70 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	69 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	87 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_1666/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(72) & convTransposeB_CP_4179_elements(70) & convTransposeB_CP_4179_elements(71) & convTransposeB_CP_4179_elements(69);
      gj_convTransposeB_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	1 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1813/SplitProtocol/Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1813/SplitProtocol/Sample/ra
      -- 
    ra_4859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1813_inst_ack_0, ack => convTransposeB_CP_4179_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	1 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1813/SplitProtocol/Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1813/SplitProtocol/Update/ca
      -- 
    ca_4864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1813_inst_ack_1, ack => convTransposeB_CP_4179_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	86 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1810/$exit
      -- CP-element group 76: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1813/$exit
      -- CP-element group 76: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_sources/type_cast_1813/SplitProtocol/$exit
      -- CP-element group 76: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1810/phi_stmt_1810_req
      -- 
    phi_stmt_1810_req_4865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1810_req_4865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(76), ack => phi_stmt_1810_req_0); -- 
    convTransposeB_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(74) & convTransposeB_CP_4179_elements(75);
      gj_convTransposeB_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	1 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/Sample/ra
      -- 
    ra_4882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1809_inst_ack_0, ack => convTransposeB_CP_4179_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	1 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/Update/ca
      -- 
    ca_4887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1809_inst_ack_1, ack => convTransposeB_CP_4179_elements(78)); -- 
    -- CP-element group 79:  join  transition  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	86 
    -- CP-element group 79:  members (5) 
      -- CP-element group 79: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1803/$exit
      -- CP-element group 79: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/$exit
      -- CP-element group 79: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_sources/type_cast_1809/SplitProtocol/$exit
      -- CP-element group 79: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1803/phi_stmt_1803_req
      -- 
    phi_stmt_1803_req_4888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1803_req_4888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(79), ack => phi_stmt_1803_req_1); -- 
    convTransposeB_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(77) & convTransposeB_CP_4179_elements(78);
      gj_convTransposeB_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	1 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/Sample/ra
      -- 
    ra_4905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1799_inst_ack_0, ack => convTransposeB_CP_4179_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	1 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/Update/ca
      -- 
    ca_4910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1799_inst_ack_1, ack => convTransposeB_CP_4179_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	86 
    -- CP-element group 82:  members (5) 
      -- CP-element group 82: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1796/$exit
      -- CP-element group 82: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/$exit
      -- CP-element group 82: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_sources/type_cast_1799/SplitProtocol/$exit
      -- CP-element group 82: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1796/phi_stmt_1796_req
      -- 
    phi_stmt_1796_req_4911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1796_req_4911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(82), ack => phi_stmt_1796_req_0); -- 
    convTransposeB_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(80) & convTransposeB_CP_4179_elements(81);
      gj_convTransposeB_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	1 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_sources/type_cast_1792/SplitProtocol/Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_sources/type_cast_1792/SplitProtocol/Sample/ra
      -- 
    ra_4928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1792_inst_ack_0, ack => convTransposeB_CP_4179_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	1 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_sources/type_cast_1792/SplitProtocol/Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_sources/type_cast_1792/SplitProtocol/Update/ca
      -- 
    ca_4933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1792_inst_ack_1, ack => convTransposeB_CP_4179_elements(84)); -- 
    -- CP-element group 85:  join  transition  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1789/$exit
      -- CP-element group 85: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_sources/$exit
      -- CP-element group 85: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_sources/type_cast_1792/$exit
      -- CP-element group 85: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_sources/type_cast_1792/SplitProtocol/$exit
      -- CP-element group 85: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/phi_stmt_1789/phi_stmt_1789_req
      -- 
    phi_stmt_1789_req_4934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1789_req_4934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(85), ack => phi_stmt_1789_req_0); -- 
    convTransposeB_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(83) & convTransposeB_CP_4179_elements(84);
      gj_convTransposeB_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  join  transition  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	76 
    -- CP-element group 86: 	79 
    -- CP-element group 86: 	82 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_1666/ifx_xend134_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(76) & convTransposeB_CP_4179_elements(79) & convTransposeB_CP_4179_elements(82) & convTransposeB_CP_4179_elements(85);
      gj_convTransposeB_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  merge  fork  transition  place  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	73 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	89 
    -- CP-element group 87: 	90 
    -- CP-element group 87: 	91 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1666/merge_stmt_1788_PhiReqMerge
      -- CP-element group 87: 	 branch_block_stmt_1666/merge_stmt_1788_PhiAck/$entry
      -- 
    convTransposeB_CP_4179_elements(87) <= OrReduce(convTransposeB_CP_4179_elements(73) & convTransposeB_CP_4179_elements(86));
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	92 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_1666/merge_stmt_1788_PhiAck/phi_stmt_1789_ack
      -- 
    phi_stmt_1789_ack_4939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1789_ack_0, ack => convTransposeB_CP_4179_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	92 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_1666/merge_stmt_1788_PhiAck/phi_stmt_1796_ack
      -- 
    phi_stmt_1796_ack_4940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1796_ack_0, ack => convTransposeB_CP_4179_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_1666/merge_stmt_1788_PhiAck/phi_stmt_1803_ack
      -- 
    phi_stmt_1803_ack_4941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1803_ack_0, ack => convTransposeB_CP_4179_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	87 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_1666/merge_stmt_1788_PhiAck/phi_stmt_1810_ack
      -- 
    phi_stmt_1810_ack_4942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1810_ack_0, ack => convTransposeB_CP_4179_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  place  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	88 
    -- CP-element group 92: 	89 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	30 
    -- CP-element group 92: 	31 
    -- CP-element group 92: 	34 
    -- CP-element group 92: 	35 
    -- CP-element group 92: 	36 
    -- CP-element group 92: 	50 
    -- CP-element group 92: 	33 
    -- CP-element group 92: 	43 
    -- CP-element group 92: 	41 
    -- CP-element group 92: 	48 
    -- CP-element group 92: 	32 
    -- CP-element group 92: 	46 
    -- CP-element group 92: 	39 
    -- CP-element group 92: 	37 
    -- CP-element group 92: 	53 
    -- CP-element group 92:  members (53) 
      -- CP-element group 92: 	 branch_block_stmt_1666/merge_stmt_1788__exit__
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944__entry__
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1830_update_start_
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1830_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1907_update_start_
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1900_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1900_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1900_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1900_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1900_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1900_update_start_
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1858_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1858_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1858_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_final_index_sum_regn_update_start
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1830_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1830_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_final_index_sum_regn_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1906_final_index_sum_regn_Update/req
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1830_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1830_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1844_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1844_update_start_
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1858_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1858_update_start_
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1844_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1844_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1844_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1844_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_update_start_
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1858_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1907_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1907_complete/req
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Update/word_access_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1911_Update/word_access_complete/word_0/cr
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1921_update_start_
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1921_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/type_cast_1921_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1928_update_start_
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_final_index_sum_regn_update_start
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_final_index_sum_regn_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/array_obj_ref_1927_final_index_sum_regn_Update/req
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1928_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/addr_of_1928_complete/req
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_update_start_
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Update/word_access_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_1666/assign_stmt_1822_to_assign_stmt_1944/ptr_deref_1931_Update/word_access_complete/word_0/cr
      -- CP-element group 92: 	 branch_block_stmt_1666/merge_stmt_1788_PhiAck/$exit
      -- 
    cr_4476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(92), ack => type_cast_1900_inst_req_1); -- 
    rr_4471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(92), ack => type_cast_1900_inst_req_0); -- 
    cr_4462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(92), ack => type_cast_1858_inst_req_1); -- 
    rr_4457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(92), ack => type_cast_1858_inst_req_0); -- 
    cr_4434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(92), ack => type_cast_1830_inst_req_1); -- 
    req_4507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(92), ack => array_obj_ref_1906_index_offset_req_1); -- 
    rr_4429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(92), ack => type_cast_1830_inst_req_0); -- 
    rr_4443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(92), ack => type_cast_1844_inst_req_0); -- 
    cr_4448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(92), ack => type_cast_1844_inst_req_1); -- 
    req_4522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(92), ack => addr_of_1907_final_reg_req_1); -- 
    cr_4567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(92), ack => ptr_deref_1911_load_0_req_1); -- 
    cr_4586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(92), ack => type_cast_1921_inst_req_1); -- 
    req_4617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(92), ack => array_obj_ref_1927_index_offset_req_1); -- 
    req_4632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(92), ack => addr_of_1928_final_reg_req_1); -- 
    cr_4682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(92), ack => ptr_deref_1931_store_0_req_1); -- 
    convTransposeB_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(88) & convTransposeB_CP_4179_elements(89) & convTransposeB_CP_4179_elements(90) & convTransposeB_CP_4179_elements(91);
      gj_convTransposeB_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	64 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2023/SplitProtocol/Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2023/SplitProtocol/Sample/ra
      -- 
    ra_4986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2023_inst_ack_0, ack => convTransposeB_CP_4179_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	64 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2023/SplitProtocol/Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2023/SplitProtocol/Update/ca
      -- 
    ca_4991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2023_inst_ack_1, ack => convTransposeB_CP_4179_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	100 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2020/$exit
      -- CP-element group 95: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2023/$exit
      -- CP-element group 95: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2023/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_req
      -- 
    phi_stmt_2020_req_4992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2020_req_4992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(95), ack => phi_stmt_2020_req_0); -- 
    convTransposeB_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(93) & convTransposeB_CP_4179_elements(94);
      gj_convTransposeB_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	64 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/Sample/ra
      -- 
    ra_5009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2017_inst_ack_0, ack => convTransposeB_CP_4179_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	64 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/Update/ca
      -- 
    ca_5014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2017_inst_ack_1, ack => convTransposeB_CP_4179_elements(97)); -- 
    -- CP-element group 98:  join  transition  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (5) 
      -- CP-element group 98: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2014/$exit
      -- CP-element group 98: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/$exit
      -- CP-element group 98: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/$exit
      -- CP-element group 98: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2017/SplitProtocol/$exit
      -- CP-element group 98: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_req
      -- 
    phi_stmt_2014_req_5015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2014_req_5015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(98), ack => phi_stmt_2014_req_0); -- 
    convTransposeB_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(96) & convTransposeB_CP_4179_elements(97);
      gj_convTransposeB_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  transition  output  delay-element  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	64 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (4) 
      -- CP-element group 99: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2007/$exit
      -- CP-element group 99: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_sources/$exit
      -- CP-element group 99: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_sources/type_cast_2011_konst_delay_trans
      -- CP-element group 99: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_req
      -- 
    phi_stmt_2007_req_5023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2007_req_5023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(99), ack => phi_stmt_2007_req_0); -- 
    -- Element group convTransposeB_CP_4179_elements(99) is a control-delay.
    cp_element_99_delay: control_delay_element  generic map(name => " 99_delay", delay_value => 1)  port map(req => convTransposeB_CP_4179_elements(64), ack => convTransposeB_CP_4179_elements(99), clk => clk, reset =>reset);
    -- CP-element group 100:  join  transition  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	95 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	111 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1666/ifx_xelse_ifx_xend134_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(95) & convTransposeB_CP_4179_elements(98) & convTransposeB_CP_4179_elements(99);
      gj_convTransposeB_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	55 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2025/SplitProtocol/Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2025/SplitProtocol/Sample/ra
      -- 
    ra_5043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2025_inst_ack_0, ack => convTransposeB_CP_4179_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	55 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2025/SplitProtocol/Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2025/SplitProtocol/Update/ca
      -- 
    ca_5048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2025_inst_ack_1, ack => convTransposeB_CP_4179_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	110 
    -- CP-element group 103:  members (5) 
      -- CP-element group 103: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2020/$exit
      -- CP-element group 103: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/$exit
      -- CP-element group 103: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2025/$exit
      -- CP-element group 103: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_sources/type_cast_2025/SplitProtocol/$exit
      -- CP-element group 103: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2020/phi_stmt_2020_req
      -- 
    phi_stmt_2020_req_5049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2020_req_5049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(103), ack => phi_stmt_2020_req_1); -- 
    convTransposeB_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(101) & convTransposeB_CP_4179_elements(102);
      gj_convTransposeB_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	55 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2019/SplitProtocol/Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2019/SplitProtocol/Sample/ra
      -- 
    ra_5066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2019_inst_ack_0, ack => convTransposeB_CP_4179_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	55 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2019/SplitProtocol/Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2019/SplitProtocol/Update/ca
      -- 
    ca_5071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2019_inst_ack_1, ack => convTransposeB_CP_4179_elements(105)); -- 
    -- CP-element group 106:  join  transition  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	110 
    -- CP-element group 106:  members (5) 
      -- CP-element group 106: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2014/$exit
      -- CP-element group 106: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/$exit
      -- CP-element group 106: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2019/$exit
      -- CP-element group 106: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_sources/type_cast_2019/SplitProtocol/$exit
      -- CP-element group 106: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2014/phi_stmt_2014_req
      -- 
    phi_stmt_2014_req_5072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2014_req_5072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(106), ack => phi_stmt_2014_req_1); -- 
    convTransposeB_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(104) & convTransposeB_CP_4179_elements(105);
      gj_convTransposeB_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	55 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_sources/type_cast_2013/SplitProtocol/Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_sources/type_cast_2013/SplitProtocol/Sample/ra
      -- 
    ra_5089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2013_inst_ack_0, ack => convTransposeB_CP_4179_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	55 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_sources/type_cast_2013/SplitProtocol/Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_sources/type_cast_2013/SplitProtocol/Update/ca
      -- 
    ca_5094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2013_inst_ack_1, ack => convTransposeB_CP_4179_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2007/$exit
      -- CP-element group 109: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_sources/$exit
      -- CP-element group 109: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_sources/type_cast_2013/$exit
      -- CP-element group 109: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_sources/type_cast_2013/SplitProtocol/$exit
      -- CP-element group 109: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/phi_stmt_2007/phi_stmt_2007_req
      -- 
    phi_stmt_2007_req_5095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2007_req_5095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_4179_elements(109), ack => phi_stmt_2007_req_1); -- 
    convTransposeB_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(107) & convTransposeB_CP_4179_elements(108);
      gj_convTransposeB_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  transition  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	103 
    -- CP-element group 110: 	106 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1666/ifx_xthen_ifx_xend134_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(103) & convTransposeB_CP_4179_elements(106) & convTransposeB_CP_4179_elements(109);
      gj_convTransposeB_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  merge  fork  transition  place  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	100 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	113 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_1666/merge_stmt_2006_PhiReqMerge
      -- CP-element group 111: 	 branch_block_stmt_1666/merge_stmt_2006_PhiAck/$entry
      -- 
    convTransposeB_CP_4179_elements(111) <= OrReduce(convTransposeB_CP_4179_elements(100) & convTransposeB_CP_4179_elements(110));
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	115 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_1666/merge_stmt_2006_PhiAck/phi_stmt_2007_ack
      -- 
    phi_stmt_2007_ack_5100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2007_ack_0, ack => convTransposeB_CP_4179_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_1666/merge_stmt_2006_PhiAck/phi_stmt_2014_ack
      -- 
    phi_stmt_2014_ack_5101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2014_ack_0, ack => convTransposeB_CP_4179_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_1666/merge_stmt_2006_PhiAck/phi_stmt_2020_ack
      -- 
    phi_stmt_2020_ack_5102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2020_ack_0, ack => convTransposeB_CP_4179_elements(114)); -- 
    -- CP-element group 115:  join  transition  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	112 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	1 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_1666/merge_stmt_2006_PhiAck/$exit
      -- 
    convTransposeB_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeB_CP_4179_elements(112) & convTransposeB_CP_4179_elements(113) & convTransposeB_CP_4179_elements(114);
      gj_convTransposeB_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_4179_elements(115), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom92_1926_resized : std_logic_vector(13 downto 0);
    signal R_idxprom92_1926_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1905_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1905_scaled : std_logic_vector(13 downto 0);
    signal add104_1957 : std_logic_vector(15 downto 0);
    signal add64_1745 : std_logic_vector(31 downto 0);
    signal add83_1881 : std_logic_vector(31 downto 0);
    signal add85_1891 : std_logic_vector(31 downto 0);
    signal add97_1939 : std_logic_vector(31 downto 0);
    signal add_1734 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_1827 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1906_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1906_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1906_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1906_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1906_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1906_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1927_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1927_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1927_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1927_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1927_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1927_root_address : std_logic_vector(13 downto 0);
    signal arrayidx88_1908 : std_logic_vector(31 downto 0);
    signal arrayidx93_1929 : std_logic_vector(31 downto 0);
    signal call10_1681 : std_logic_vector(31 downto 0);
    signal call13_1684 : std_logic_vector(31 downto 0);
    signal call16_1687 : std_logic_vector(31 downto 0);
    signal call19_1690 : std_logic_vector(31 downto 0);
    signal call1_1672 : std_logic_vector(31 downto 0);
    signal call21_1693 : std_logic_vector(31 downto 0);
    signal call23_1696 : std_logic_vector(31 downto 0);
    signal call24_1699 : std_logic_vector(31 downto 0);
    signal call27_1702 : std_logic_vector(31 downto 0);
    signal call30_1705 : std_logic_vector(31 downto 0);
    signal call4_1675 : std_logic_vector(31 downto 0);
    signal call7_1678 : std_logic_vector(31 downto 0);
    signal call_1669 : std_logic_vector(31 downto 0);
    signal cmp112_1974 : std_logic_vector(0 downto 0);
    signal cmp123_1999 : std_logic_vector(0 downto 0);
    signal cmp_1944 : std_logic_vector(0 downto 0);
    signal conv100_1768 : std_logic_vector(31 downto 0);
    signal conv108_1969 : std_logic_vector(31 downto 0);
    signal conv111_1774 : std_logic_vector(31 downto 0);
    signal conv118_1994 : std_logic_vector(31 downto 0);
    signal conv121_1780 : std_logic_vector(31 downto 0);
    signal conv34_1712 : std_logic_vector(31 downto 0);
    signal conv35_1722 : std_logic_vector(15 downto 0);
    signal conv46_1831 : std_logic_vector(31 downto 0);
    signal conv48_1728 : std_logic_vector(31 downto 0);
    signal conv57_1845 : std_logic_vector(31 downto 0);
    signal conv71_1859 : std_logic_vector(31 downto 0);
    signal conv74_1756 : std_logic_vector(31 downto 0);
    signal conv76_1865 : std_logic_vector(31 downto 0);
    signal conv79_1762 : std_logic_vector(31 downto 0);
    signal conv81_1871 : std_logic_vector(31 downto 0);
    signal idxprom92_1922 : std_logic_vector(63 downto 0);
    signal idxprom_1901 : std_logic_vector(63 downto 0);
    signal inc116_1978 : std_logic_vector(15 downto 0);
    signal inc116x_xinput_dim0x_x2_1983 : std_logic_vector(15 downto 0);
    signal inc_1965 : std_logic_vector(15 downto 0);
    signal indvar_1789 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2032 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2020 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_1810 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2014 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_1803 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1990 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2007 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1796 : std_logic_vector(15 downto 0);
    signal mul60_1850 : std_logic_vector(31 downto 0);
    signal mul82_1876 : std_logic_vector(31 downto 0);
    signal mul84_1886 : std_logic_vector(31 downto 0);
    signal mul_1836 : std_logic_vector(31 downto 0);
    signal ptr_deref_1911_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1911_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1911_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1911_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1911_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1931_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1931_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1931_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1931_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1931_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1931_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr122138_1786 : std_logic_vector(31 downto 0);
    signal shr137_1718 : std_logic_vector(31 downto 0);
    signal shr87_1897 : std_logic_vector(31 downto 0);
    signal shr91_1918 : std_logic_vector(31 downto 0);
    signal sub54_1841 : std_logic_vector(31 downto 0);
    signal sub67_1750 : std_logic_vector(31 downto 0);
    signal sub68_1855 : std_logic_vector(31 downto 0);
    signal sub_1739 : std_logic_vector(31 downto 0);
    signal tmp1_1822 : std_logic_vector(31 downto 0);
    signal tmp89_1912 : std_logic_vector(63 downto 0);
    signal type_cast_1710_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1716_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1726_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1732_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1743_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1754_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1760_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1766_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1772_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1778_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1784_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1792_wire : std_logic_vector(31 downto 0);
    signal type_cast_1795_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1799_wire : std_logic_vector(15 downto 0);
    signal type_cast_1802_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1807_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1809_wire : std_logic_vector(15 downto 0);
    signal type_cast_1813_wire : std_logic_vector(15 downto 0);
    signal type_cast_1815_wire : std_logic_vector(15 downto 0);
    signal type_cast_1820_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1863_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1869_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1895_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1916_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1937_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1955_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1963_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1987_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2011_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2013_wire : std_logic_vector(15 downto 0);
    signal type_cast_2017_wire : std_logic_vector(15 downto 0);
    signal type_cast_2019_wire : std_logic_vector(15 downto 0);
    signal type_cast_2023_wire : std_logic_vector(15 downto 0);
    signal type_cast_2025_wire : std_logic_vector(15 downto 0);
    signal type_cast_2030_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2038_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1906_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1906_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1906_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1906_resized_base_address <= "00000000000000";
    array_obj_ref_1927_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1927_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1927_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1927_resized_base_address <= "00000000000000";
    ptr_deref_1911_word_offset_0 <= "00000000000000";
    ptr_deref_1931_word_offset_0 <= "00000000000000";
    type_cast_1710_wire_constant <= "00000000000000000000000000000010";
    type_cast_1716_wire_constant <= "00000000000000000011111111111111";
    type_cast_1726_wire_constant <= "00000000000000001111111111111111";
    type_cast_1732_wire_constant <= "00000000000000001111111111111111";
    type_cast_1743_wire_constant <= "00000000000000001111111111111111";
    type_cast_1754_wire_constant <= "00000000000000001111111111111111";
    type_cast_1760_wire_constant <= "00000000000000001111111111111111";
    type_cast_1766_wire_constant <= "00000000000000001111111111111111";
    type_cast_1772_wire_constant <= "00000000000000001111111111111111";
    type_cast_1778_wire_constant <= "00000000000000000000000000000001";
    type_cast_1784_wire_constant <= "00000000000000000111111111111111";
    type_cast_1795_wire_constant <= "00000000000000000000000000000000";
    type_cast_1802_wire_constant <= "0000000000000000";
    type_cast_1807_wire_constant <= "0000000000000000";
    type_cast_1820_wire_constant <= "00000000000000000000000000000100";
    type_cast_1863_wire_constant <= "00000000000000001111111111111111";
    type_cast_1869_wire_constant <= "00000000000000001111111111111111";
    type_cast_1895_wire_constant <= "00000000000000000000000000000010";
    type_cast_1916_wire_constant <= "00000000000000000000000000000010";
    type_cast_1937_wire_constant <= "00000000000000000000000000000100";
    type_cast_1955_wire_constant <= "0000000000000100";
    type_cast_1963_wire_constant <= "0000000000000001";
    type_cast_1987_wire_constant <= "0000000000000000";
    type_cast_2011_wire_constant <= "0000000000000000";
    type_cast_2030_wire_constant <= "00000000000000000000000000000001";
    type_cast_2038_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_1789: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1792_wire & type_cast_1795_wire_constant;
      req <= phi_stmt_1789_req_0 & phi_stmt_1789_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1789",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1789_ack_0,
          idata => idata,
          odata => indvar_1789,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1789
    phi_stmt_1796: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1799_wire & type_cast_1802_wire_constant;
      req <= phi_stmt_1796_req_0 & phi_stmt_1796_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1796",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1796_ack_0,
          idata => idata,
          odata => input_dim2x_x1_1796,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1796
    phi_stmt_1803: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1807_wire_constant & type_cast_1809_wire;
      req <= phi_stmt_1803_req_0 & phi_stmt_1803_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1803",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1803_ack_0,
          idata => idata,
          odata => input_dim1x_x1_1803,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1803
    phi_stmt_1810: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1813_wire & type_cast_1815_wire;
      req <= phi_stmt_1810_req_0 & phi_stmt_1810_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1810",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1810_ack_0,
          idata => idata,
          odata => input_dim0x_x2_1810,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1810
    phi_stmt_2007: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2011_wire_constant & type_cast_2013_wire;
      req <= phi_stmt_2007_req_0 & phi_stmt_2007_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2007",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2007_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2007,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2007
    phi_stmt_2014: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2017_wire & type_cast_2019_wire;
      req <= phi_stmt_2014_req_0 & phi_stmt_2014_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2014",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2014_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2014,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2014
    phi_stmt_2020: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2023_wire & type_cast_2025_wire;
      req <= phi_stmt_2020_req_0 & phi_stmt_2020_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2020",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2020_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2020,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2020
    -- flow-through select operator MUX_1989_inst
    input_dim1x_x2_1990 <= type_cast_1987_wire_constant when (cmp112_1974(0) /=  '0') else inc_1965;
    addr_of_1907_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1907_final_reg_req_0;
      addr_of_1907_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1907_final_reg_req_1;
      addr_of_1907_final_reg_ack_1<= rack(0);
      addr_of_1907_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1907_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1906_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx88_1908,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1928_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1928_final_reg_req_0;
      addr_of_1928_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1928_final_reg_req_1;
      addr_of_1928_final_reg_ack_1<= rack(0);
      addr_of_1928_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1928_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1927_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx93_1929,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1721_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1721_inst_req_0;
      type_cast_1721_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1721_inst_req_1;
      type_cast_1721_inst_ack_1<= rack(0);
      type_cast_1721_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1721_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr137_1718,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_1722,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1792_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1792_inst_req_0;
      type_cast_1792_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1792_inst_req_1;
      type_cast_1792_inst_ack_1<= rack(0);
      type_cast_1792_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1792_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2032,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1792_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1799_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1799_inst_req_0;
      type_cast_1799_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1799_inst_req_1;
      type_cast_1799_inst_ack_1<= rack(0);
      type_cast_1799_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1799_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2007,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1799_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1809_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1809_inst_req_0;
      type_cast_1809_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1809_inst_req_1;
      type_cast_1809_inst_ack_1<= rack(0);
      type_cast_1809_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1809_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2014,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1809_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1813_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1813_inst_req_0;
      type_cast_1813_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1813_inst_req_1;
      type_cast_1813_inst_ack_1<= rack(0);
      type_cast_1813_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1813_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2020,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1813_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1815_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1815_inst_req_0;
      type_cast_1815_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1815_inst_req_1;
      type_cast_1815_inst_ack_1<= rack(0);
      type_cast_1815_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1815_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv35_1722,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1815_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1830_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1830_inst_req_0;
      type_cast_1830_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1830_inst_req_1;
      type_cast_1830_inst_ack_1<= rack(0);
      type_cast_1830_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1830_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1810,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv46_1831,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1844_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1844_inst_req_0;
      type_cast_1844_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1844_inst_req_1;
      type_cast_1844_inst_ack_1<= rack(0);
      type_cast_1844_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1844_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1803,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv57_1845,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1858_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1858_inst_req_0;
      type_cast_1858_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1858_inst_req_1;
      type_cast_1858_inst_ack_1<= rack(0);
      type_cast_1858_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1858_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1796,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_1859,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1900_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1900_inst_req_0;
      type_cast_1900_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1900_inst_req_1;
      type_cast_1900_inst_ack_1<= rack(0);
      type_cast_1900_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1900_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr87_1897,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1901,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1921_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1921_inst_req_0;
      type_cast_1921_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1921_inst_req_1;
      type_cast_1921_inst_ack_1<= rack(0);
      type_cast_1921_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1921_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr91_1918,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom92_1922,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1968_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1968_inst_req_0;
      type_cast_1968_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1968_inst_req_1;
      type_cast_1968_inst_ack_1<= rack(0);
      type_cast_1968_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1968_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_1965,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv108_1969,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1977_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1977_inst_req_0;
      type_cast_1977_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1977_inst_req_1;
      type_cast_1977_inst_ack_1<= rack(0);
      type_cast_1977_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1977_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp112_1974,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc116_1978,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1993_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1993_inst_req_0;
      type_cast_1993_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1993_inst_req_1;
      type_cast_1993_inst_ack_1<= rack(0);
      type_cast_1993_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1993_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc116x_xinput_dim0x_x2_1983,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv118_1994,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2013_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2013_inst_req_0;
      type_cast_2013_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2013_inst_req_1;
      type_cast_2013_inst_ack_1<= rack(0);
      type_cast_2013_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2013_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add104_1957,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2013_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2017_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2017_inst_req_0;
      type_cast_2017_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2017_inst_req_1;
      type_cast_2017_inst_ack_1<= rack(0);
      type_cast_2017_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2017_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1990,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2017_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2019_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2019_inst_req_0;
      type_cast_2019_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2019_inst_req_1;
      type_cast_2019_inst_ack_1<= rack(0);
      type_cast_2019_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2019_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_1803,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2019_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2023_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2023_inst_req_0;
      type_cast_2023_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2023_inst_req_1;
      type_cast_2023_inst_ack_1<= rack(0);
      type_cast_2023_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2023_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc116x_xinput_dim0x_x2_1983,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2023_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2025_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2025_inst_req_0;
      type_cast_2025_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2025_inst_req_1;
      type_cast_2025_inst_ack_1<= rack(0);
      type_cast_2025_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2025_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_1810,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2025_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1906_index_1_rename
    process(R_idxprom_1905_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1905_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1905_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1906_index_1_resize
    process(idxprom_1901) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1901;
      ov := iv(13 downto 0);
      R_idxprom_1905_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1906_root_address_inst
    process(array_obj_ref_1906_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1906_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1906_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1927_index_1_rename
    process(R_idxprom92_1926_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom92_1926_resized;
      ov(13 downto 0) := iv;
      R_idxprom92_1926_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1927_index_1_resize
    process(idxprom92_1922) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom92_1922;
      ov := iv(13 downto 0);
      R_idxprom92_1926_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1927_root_address_inst
    process(array_obj_ref_1927_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1927_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1927_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1911_addr_0
    process(ptr_deref_1911_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1911_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1911_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1911_base_resize
    process(arrayidx88_1908) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx88_1908;
      ov := iv(13 downto 0);
      ptr_deref_1911_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1911_gather_scatter
    process(ptr_deref_1911_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1911_data_0;
      ov(63 downto 0) := iv;
      tmp89_1912 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1911_root_address_inst
    process(ptr_deref_1911_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1911_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1911_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1931_addr_0
    process(ptr_deref_1931_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1931_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1931_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1931_base_resize
    process(arrayidx93_1929) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx93_1929;
      ov := iv(13 downto 0);
      ptr_deref_1931_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1931_gather_scatter
    process(tmp89_1912) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp89_1912;
      ov(63 downto 0) := iv;
      ptr_deref_1931_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1931_root_address_inst
    process(ptr_deref_1931_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1931_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1931_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1945_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1944;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1945_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1945_branch_req_0,
          ack0 => if_stmt_1945_branch_ack_0,
          ack1 => if_stmt_1945_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2000_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp123_1999;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2000_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2000_branch_req_0,
          ack0 => if_stmt_2000_branch_ack_0,
          ack1 => if_stmt_2000_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1956_inst
    process(input_dim2x_x1_1796) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_1796, type_cast_1955_wire_constant, tmp_var);
      add104_1957 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1964_inst
    process(input_dim1x_x1_1803) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_1803, type_cast_1963_wire_constant, tmp_var);
      inc_1965 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1982_inst
    process(inc116_1978, input_dim0x_x2_1810) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc116_1978, input_dim0x_x2_1810, tmp_var);
      inc116x_xinput_dim0x_x2_1983 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1733_inst
    process(call10_1681) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call10_1681, type_cast_1732_wire_constant, tmp_var);
      add_1734 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1744_inst
    process(call13_1684) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call13_1684, type_cast_1743_wire_constant, tmp_var);
      add64_1745 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1826_inst
    process(call23_1696, tmp1_1822) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call23_1696, tmp1_1822, tmp_var);
      add_src_0x_x0_1827 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1840_inst
    process(sub_1739, mul_1836) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_1739, mul_1836, tmp_var);
      sub54_1841 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1854_inst
    process(sub67_1750, mul60_1850) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub67_1750, mul60_1850, tmp_var);
      sub68_1855 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1880_inst
    process(mul82_1876, conv76_1865) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul82_1876, conv76_1865, tmp_var);
      add83_1881 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1890_inst
    process(mul84_1886, conv71_1859) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul84_1886, conv71_1859, tmp_var);
      add85_1891 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1938_inst
    process(conv71_1859) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv71_1859, type_cast_1937_wire_constant, tmp_var);
      add97_1939 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2031_inst
    process(indvar_1789) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1789, type_cast_2030_wire_constant, tmp_var);
      indvarx_xnext_2032 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1717_inst
    process(conv34_1712) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv34_1712, type_cast_1716_wire_constant, tmp_var);
      shr137_1718 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1727_inst
    process(call19_1690) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call19_1690, type_cast_1726_wire_constant, tmp_var);
      conv48_1728 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1755_inst
    process(call30_1705) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call30_1705, type_cast_1754_wire_constant, tmp_var);
      conv74_1756 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1761_inst
    process(call27_1702) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call27_1702, type_cast_1760_wire_constant, tmp_var);
      conv79_1762 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1767_inst
    process(call4_1675) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call4_1675, type_cast_1766_wire_constant, tmp_var);
      conv100_1768 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1773_inst
    process(call1_1672) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call1_1672, type_cast_1772_wire_constant, tmp_var);
      conv111_1774 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1785_inst
    process(conv121_1780) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv121_1780, type_cast_1784_wire_constant, tmp_var);
      shr122138_1786 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1864_inst
    process(sub68_1855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(sub68_1855, type_cast_1863_wire_constant, tmp_var);
      conv76_1865 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1870_inst
    process(sub54_1841) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(sub54_1841, type_cast_1869_wire_constant, tmp_var);
      conv81_1871 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1973_inst
    process(conv108_1969, conv111_1774) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv108_1969, conv111_1774, tmp_var);
      cmp112_1974 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1998_inst
    process(conv118_1994, shr122138_1786) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv118_1994, shr122138_1786, tmp_var);
      cmp123_1999 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1711_inst
    process(call_1669) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1669, type_cast_1710_wire_constant, tmp_var);
      conv34_1712 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1779_inst
    process(call_1669) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_1669, type_cast_1778_wire_constant, tmp_var);
      conv121_1780 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1896_inst
    process(add_src_0x_x0_1827) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_1827, type_cast_1895_wire_constant, tmp_var);
      shr87_1897 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1917_inst
    process(add85_1891) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add85_1891, type_cast_1916_wire_constant, tmp_var);
      shr91_1918 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1821_inst
    process(indvar_1789) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1789, type_cast_1820_wire_constant, tmp_var);
      tmp1_1822 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1835_inst
    process(conv46_1831, conv48_1728) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv46_1831, conv48_1728, tmp_var);
      mul_1836 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1849_inst
    process(conv57_1845, conv48_1728) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv57_1845, conv48_1728, tmp_var);
      mul60_1850 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1875_inst
    process(conv81_1871, conv79_1762) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv81_1871, conv79_1762, tmp_var);
      mul82_1876 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1885_inst
    process(add83_1881, conv74_1756) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add83_1881, conv74_1756, tmp_var);
      mul84_1886 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1738_inst
    process(add_1734, call21_1693) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add_1734, call21_1693, tmp_var);
      sub_1739 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1749_inst
    process(add64_1745, call21_1693) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add64_1745, call21_1693, tmp_var);
      sub67_1750 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1943_inst
    process(add97_1939, conv100_1768) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add97_1939, conv100_1768, tmp_var);
      cmp_1944 <= tmp_var; --
    end process;
    -- shared split operator group (35) : array_obj_ref_1906_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1905_scaled;
      array_obj_ref_1906_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1906_index_offset_req_0;
      array_obj_ref_1906_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1906_index_offset_req_1;
      array_obj_ref_1906_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : array_obj_ref_1927_index_offset 
    ApIntAdd_group_36: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom92_1926_scaled;
      array_obj_ref_1927_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1927_index_offset_req_0;
      array_obj_ref_1927_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1927_index_offset_req_1;
      array_obj_ref_1927_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_36_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared load operator group (0) : ptr_deref_1911_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1911_load_0_req_0;
      ptr_deref_1911_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1911_load_0_req_1;
      ptr_deref_1911_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1911_word_address_0;
      ptr_deref_1911_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1931_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1931_store_0_req_0;
      ptr_deref_1931_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1931_store_0_req_1;
      ptr_deref_1931_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1931_word_address_0;
      data_in <= ptr_deref_1931_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1668_inst RPIPE_Block1_start_1671_inst RPIPE_Block1_start_1674_inst RPIPE_Block1_start_1677_inst RPIPE_Block1_start_1680_inst RPIPE_Block1_start_1683_inst RPIPE_Block1_start_1686_inst RPIPE_Block1_start_1689_inst RPIPE_Block1_start_1692_inst RPIPE_Block1_start_1695_inst RPIPE_Block1_start_1698_inst RPIPE_Block1_start_1701_inst RPIPE_Block1_start_1704_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(415 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 12 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 12 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 12 downto 0);
      signal guard_vector : std_logic_vector( 12 downto 0);
      constant outBUFs : IntegerArray(12 downto 0) := (12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(12 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false);
      constant guardBuffering: IntegerArray(12 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2);
      -- 
    begin -- 
      reqL_unguarded(12) <= RPIPE_Block1_start_1668_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block1_start_1671_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block1_start_1674_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block1_start_1677_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block1_start_1680_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block1_start_1683_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block1_start_1686_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block1_start_1689_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block1_start_1692_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block1_start_1695_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block1_start_1698_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block1_start_1701_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block1_start_1704_inst_req_0;
      RPIPE_Block1_start_1668_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block1_start_1671_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block1_start_1674_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block1_start_1677_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block1_start_1680_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block1_start_1683_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block1_start_1686_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block1_start_1689_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block1_start_1692_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block1_start_1695_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block1_start_1698_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block1_start_1701_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block1_start_1704_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(12) <= RPIPE_Block1_start_1668_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block1_start_1671_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block1_start_1674_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block1_start_1677_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block1_start_1680_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block1_start_1683_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block1_start_1686_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block1_start_1689_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block1_start_1692_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block1_start_1695_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block1_start_1698_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block1_start_1701_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block1_start_1704_inst_req_1;
      RPIPE_Block1_start_1668_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block1_start_1671_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block1_start_1674_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block1_start_1677_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block1_start_1680_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block1_start_1683_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block1_start_1686_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block1_start_1689_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block1_start_1692_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block1_start_1695_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block1_start_1698_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block1_start_1701_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block1_start_1704_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      call_1669 <= data_out(415 downto 384);
      call1_1672 <= data_out(383 downto 352);
      call4_1675 <= data_out(351 downto 320);
      call7_1678 <= data_out(319 downto 288);
      call10_1681 <= data_out(287 downto 256);
      call13_1684 <= data_out(255 downto 224);
      call16_1687 <= data_out(223 downto 192);
      call19_1690 <= data_out(191 downto 160);
      call21_1693 <= data_out(159 downto 128);
      call23_1696 <= data_out(127 downto 96);
      call24_1699 <= data_out(95 downto 64);
      call27_1702 <= data_out(63 downto 32);
      call30_1705 <= data_out(31 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 13, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 32,  num_reqs => 13,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2036_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2036_inst_req_0;
      WPIPE_Block1_done_2036_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2036_inst_req_1;
      WPIPE_Block1_done_2036_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2038_wire_constant;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(31 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_5119_start: Boolean;
  signal convTransposeC_CP_5119_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2100_inst_req_1 : boolean;
  signal array_obj_ref_2290_index_offset_req_0 : boolean;
  signal RPIPE_Block2_start_2077_inst_ack_1 : boolean;
  signal array_obj_ref_2290_index_offset_ack_0 : boolean;
  signal RPIPE_Block2_start_2077_inst_req_1 : boolean;
  signal array_obj_ref_2290_index_offset_req_1 : boolean;
  signal RPIPE_Block2_start_2083_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2080_inst_ack_1 : boolean;
  signal array_obj_ref_2290_index_offset_ack_1 : boolean;
  signal type_cast_2228_inst_req_0 : boolean;
  signal ptr_deref_2295_load_0_req_1 : boolean;
  signal type_cast_2100_inst_ack_1 : boolean;
  signal type_cast_2228_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2083_inst_req_1 : boolean;
  signal ptr_deref_2295_load_0_ack_1 : boolean;
  signal RPIPE_Block2_start_2083_inst_ack_1 : boolean;
  signal type_cast_2228_inst_req_1 : boolean;
  signal type_cast_2228_inst_ack_1 : boolean;
  signal type_cast_2305_inst_req_0 : boolean;
  signal addr_of_2291_final_reg_req_0 : boolean;
  signal type_cast_2305_inst_ack_0 : boolean;
  signal addr_of_2291_final_reg_ack_0 : boolean;
  signal RPIPE_Block2_start_2083_inst_req_0 : boolean;
  signal type_cast_2305_inst_req_1 : boolean;
  signal type_cast_2305_inst_ack_1 : boolean;
  signal addr_of_2291_final_reg_req_1 : boolean;
  signal RPIPE_Block2_start_2080_inst_req_0 : boolean;
  signal addr_of_2291_final_reg_ack_1 : boolean;
  signal type_cast_2242_inst_req_0 : boolean;
  signal type_cast_2242_inst_ack_0 : boolean;
  signal ptr_deref_2295_load_0_req_0 : boolean;
  signal array_obj_ref_2311_index_offset_req_0 : boolean;
  signal type_cast_2214_inst_req_0 : boolean;
  signal type_cast_2242_inst_req_1 : boolean;
  signal type_cast_2242_inst_ack_1 : boolean;
  signal type_cast_2214_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2080_inst_ack_0 : boolean;
  signal ptr_deref_2295_load_0_ack_0 : boolean;
  signal type_cast_2284_inst_req_0 : boolean;
  signal type_cast_2214_inst_req_1 : boolean;
  signal type_cast_2284_inst_ack_0 : boolean;
  signal type_cast_2214_inst_ack_1 : boolean;
  signal addr_of_2312_final_reg_req_1 : boolean;
  signal addr_of_2312_final_reg_req_0 : boolean;
  signal type_cast_2284_inst_req_1 : boolean;
  signal addr_of_2312_final_reg_ack_0 : boolean;
  signal RPIPE_Block2_start_2080_inst_req_1 : boolean;
  signal type_cast_2284_inst_ack_1 : boolean;
  signal addr_of_2312_final_reg_ack_1 : boolean;
  signal array_obj_ref_2311_index_offset_req_1 : boolean;
  signal array_obj_ref_2311_index_offset_ack_1 : boolean;
  signal type_cast_2100_inst_ack_0 : boolean;
  signal array_obj_ref_2311_index_offset_ack_0 : boolean;
  signal type_cast_2100_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2047_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2047_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2047_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2047_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2050_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2050_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2050_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2050_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2053_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2053_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2053_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2053_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2056_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2056_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2056_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2056_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2059_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2059_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2059_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2059_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2062_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2062_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2062_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2062_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2065_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2065_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2065_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2065_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2068_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2068_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2068_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2068_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2071_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2071_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2071_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2071_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2074_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2074_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2074_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2074_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2077_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2077_inst_ack_0 : boolean;
  signal ptr_deref_2315_store_0_req_0 : boolean;
  signal ptr_deref_2315_store_0_ack_0 : boolean;
  signal ptr_deref_2315_store_0_req_1 : boolean;
  signal ptr_deref_2315_store_0_ack_1 : boolean;
  signal if_stmt_2329_branch_req_0 : boolean;
  signal if_stmt_2329_branch_ack_1 : boolean;
  signal if_stmt_2329_branch_ack_0 : boolean;
  signal type_cast_2352_inst_req_0 : boolean;
  signal type_cast_2352_inst_ack_0 : boolean;
  signal type_cast_2352_inst_req_1 : boolean;
  signal type_cast_2352_inst_ack_1 : boolean;
  signal type_cast_2361_inst_req_0 : boolean;
  signal type_cast_2361_inst_ack_0 : boolean;
  signal type_cast_2361_inst_req_1 : boolean;
  signal type_cast_2361_inst_ack_1 : boolean;
  signal type_cast_2377_inst_req_0 : boolean;
  signal type_cast_2377_inst_ack_0 : boolean;
  signal type_cast_2377_inst_req_1 : boolean;
  signal type_cast_2377_inst_ack_1 : boolean;
  signal if_stmt_2384_branch_req_0 : boolean;
  signal if_stmt_2384_branch_ack_1 : boolean;
  signal if_stmt_2384_branch_ack_0 : boolean;
  signal WPIPE_Block2_done_2420_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2420_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2420_inst_req_1 : boolean;
  signal WPIPE_Block2_done_2420_inst_ack_1 : boolean;
  signal type_cast_2197_inst_req_0 : boolean;
  signal type_cast_2197_inst_ack_0 : boolean;
  signal type_cast_2197_inst_req_1 : boolean;
  signal type_cast_2197_inst_ack_1 : boolean;
  signal phi_stmt_2194_req_0 : boolean;
  signal phi_stmt_2187_req_1 : boolean;
  signal phi_stmt_2180_req_0 : boolean;
  signal phi_stmt_2173_req_0 : boolean;
  signal type_cast_2199_inst_req_0 : boolean;
  signal type_cast_2199_inst_ack_0 : boolean;
  signal type_cast_2199_inst_req_1 : boolean;
  signal type_cast_2199_inst_ack_1 : boolean;
  signal phi_stmt_2194_req_1 : boolean;
  signal type_cast_2190_inst_req_0 : boolean;
  signal type_cast_2190_inst_ack_0 : boolean;
  signal type_cast_2190_inst_req_1 : boolean;
  signal type_cast_2190_inst_ack_1 : boolean;
  signal phi_stmt_2187_req_0 : boolean;
  signal type_cast_2186_inst_req_0 : boolean;
  signal type_cast_2186_inst_ack_0 : boolean;
  signal type_cast_2186_inst_req_1 : boolean;
  signal type_cast_2186_inst_ack_1 : boolean;
  signal phi_stmt_2180_req_1 : boolean;
  signal type_cast_2179_inst_req_0 : boolean;
  signal type_cast_2179_inst_ack_0 : boolean;
  signal type_cast_2179_inst_req_1 : boolean;
  signal type_cast_2179_inst_ack_1 : boolean;
  signal phi_stmt_2173_req_1 : boolean;
  signal phi_stmt_2173_ack_0 : boolean;
  signal phi_stmt_2180_ack_0 : boolean;
  signal phi_stmt_2187_ack_0 : boolean;
  signal phi_stmt_2194_ack_0 : boolean;
  signal phi_stmt_2391_req_0 : boolean;
  signal type_cast_2401_inst_req_0 : boolean;
  signal type_cast_2401_inst_ack_0 : boolean;
  signal type_cast_2401_inst_req_1 : boolean;
  signal type_cast_2401_inst_ack_1 : boolean;
  signal phi_stmt_2398_req_0 : boolean;
  signal type_cast_2407_inst_req_0 : boolean;
  signal type_cast_2407_inst_ack_0 : boolean;
  signal type_cast_2407_inst_req_1 : boolean;
  signal type_cast_2407_inst_ack_1 : boolean;
  signal phi_stmt_2404_req_0 : boolean;
  signal type_cast_2397_inst_req_0 : boolean;
  signal type_cast_2397_inst_ack_0 : boolean;
  signal type_cast_2397_inst_req_1 : boolean;
  signal type_cast_2397_inst_ack_1 : boolean;
  signal phi_stmt_2391_req_1 : boolean;
  signal type_cast_2403_inst_req_0 : boolean;
  signal type_cast_2403_inst_ack_0 : boolean;
  signal type_cast_2403_inst_req_1 : boolean;
  signal type_cast_2403_inst_ack_1 : boolean;
  signal phi_stmt_2398_req_1 : boolean;
  signal type_cast_2409_inst_req_0 : boolean;
  signal type_cast_2409_inst_ack_0 : boolean;
  signal type_cast_2409_inst_req_1 : boolean;
  signal type_cast_2409_inst_ack_1 : boolean;
  signal phi_stmt_2404_req_1 : boolean;
  signal phi_stmt_2391_ack_0 : boolean;
  signal phi_stmt_2398_ack_0 : boolean;
  signal phi_stmt_2404_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_5119_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5119_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_5119_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_5119_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_5119: Block -- control-path 
    signal convTransposeC_CP_5119_elements: BooleanArray(115 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_5119_elements(0) <= convTransposeC_CP_5119_start;
    convTransposeC_CP_5119_symbol <= convTransposeC_CP_5119_elements(66);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2045/$entry
      -- CP-element group 0: 	 branch_block_stmt_2045/branch_block_stmt_2045__entry__
      -- CP-element group 0: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084__entry__
      -- CP-element group 0: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/$entry
      -- CP-element group 0: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2047_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2047_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2047_Sample/rr
      -- 
    rr_5167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(0), ack => RPIPE_Block2_start_2047_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	115 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	74 
    -- CP-element group 1: 	75 
    -- CP-element group 1: 	77 
    -- CP-element group 1: 	78 
    -- CP-element group 1: 	80 
    -- CP-element group 1: 	81 
    -- CP-element group 1: 	83 
    -- CP-element group 1: 	84 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2045/merge_stmt_2390__exit__
      -- CP-element group 1: 	 branch_block_stmt_2045/assign_stmt_2416__entry__
      -- CP-element group 1: 	 branch_block_stmt_2045/assign_stmt_2416__exit__
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2045/assign_stmt_2416/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/assign_stmt_2416/$exit
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2194/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2187/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2190/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2190/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2190/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2190/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2190/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2190/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2180/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_sources/type_cast_2186/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_sources/type_cast_2186/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_sources/type_cast_2186/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_sources/type_cast_2186/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_sources/type_cast_2186/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_sources/type_cast_2186/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2173/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_sources/type_cast_2179/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_sources/type_cast_2179/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_sources/type_cast_2179/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_sources/type_cast_2179/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_sources/type_cast_2179/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_sources/type_cast_2179/SplitProtocol/Update/cr
      -- 
    rr_5798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(1), ack => type_cast_2199_inst_req_0); -- 
    cr_5803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(1), ack => type_cast_2199_inst_req_1); -- 
    rr_5821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(1), ack => type_cast_2190_inst_req_0); -- 
    cr_5826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(1), ack => type_cast_2190_inst_req_1); -- 
    rr_5844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(1), ack => type_cast_2186_inst_req_0); -- 
    cr_5849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(1), ack => type_cast_2186_inst_req_1); -- 
    rr_5867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(1), ack => type_cast_2179_inst_req_0); -- 
    cr_5872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(1), ack => type_cast_2179_inst_req_1); -- 
    convTransposeC_CP_5119_elements(1) <= convTransposeC_CP_5119_elements(115);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2047_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2047_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2047_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2047_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2047_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2047_Update/cr
      -- 
    ra_5168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2047_inst_ack_0, ack => convTransposeC_CP_5119_elements(2)); -- 
    cr_5172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(2), ack => RPIPE_Block2_start_2047_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2047_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2047_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2047_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2050_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2050_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2050_Sample/rr
      -- 
    ca_5173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2047_inst_ack_1, ack => convTransposeC_CP_5119_elements(3)); -- 
    rr_5181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(3), ack => RPIPE_Block2_start_2050_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2050_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2050_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2050_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2050_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2050_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2050_Update/cr
      -- 
    ra_5182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2050_inst_ack_0, ack => convTransposeC_CP_5119_elements(4)); -- 
    cr_5186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(4), ack => RPIPE_Block2_start_2050_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2050_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2050_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2050_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2053_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2053_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2053_Sample/rr
      -- 
    ca_5187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2050_inst_ack_1, ack => convTransposeC_CP_5119_elements(5)); -- 
    rr_5195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(5), ack => RPIPE_Block2_start_2053_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2053_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2053_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2053_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2053_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2053_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2053_Update/cr
      -- 
    ra_5196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2053_inst_ack_0, ack => convTransposeC_CP_5119_elements(6)); -- 
    cr_5200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(6), ack => RPIPE_Block2_start_2053_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2053_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2053_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2053_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2056_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2056_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2056_Sample/rr
      -- 
    ca_5201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2053_inst_ack_1, ack => convTransposeC_CP_5119_elements(7)); -- 
    rr_5209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(7), ack => RPIPE_Block2_start_2056_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2056_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2056_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2056_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2056_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2056_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2056_Update/cr
      -- 
    ra_5210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2056_inst_ack_0, ack => convTransposeC_CP_5119_elements(8)); -- 
    cr_5214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(8), ack => RPIPE_Block2_start_2056_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2056_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2056_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2056_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2059_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2059_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2059_Sample/rr
      -- 
    ca_5215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2056_inst_ack_1, ack => convTransposeC_CP_5119_elements(9)); -- 
    rr_5223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(9), ack => RPIPE_Block2_start_2059_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2059_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2059_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2059_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2059_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2059_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2059_Update/cr
      -- 
    ra_5224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2059_inst_ack_0, ack => convTransposeC_CP_5119_elements(10)); -- 
    cr_5228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(10), ack => RPIPE_Block2_start_2059_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2059_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2059_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2059_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2062_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2062_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2062_Sample/rr
      -- 
    ca_5229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2059_inst_ack_1, ack => convTransposeC_CP_5119_elements(11)); -- 
    rr_5237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(11), ack => RPIPE_Block2_start_2062_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2062_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2062_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2062_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2062_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2062_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2062_Update/cr
      -- 
    ra_5238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2062_inst_ack_0, ack => convTransposeC_CP_5119_elements(12)); -- 
    cr_5242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(12), ack => RPIPE_Block2_start_2062_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2062_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2062_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2062_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2065_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2065_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2065_Sample/rr
      -- 
    ca_5243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2062_inst_ack_1, ack => convTransposeC_CP_5119_elements(13)); -- 
    rr_5251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(13), ack => RPIPE_Block2_start_2065_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2065_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2065_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2065_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2065_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2065_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2065_Update/cr
      -- 
    ra_5252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2065_inst_ack_0, ack => convTransposeC_CP_5119_elements(14)); -- 
    cr_5256_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5256_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(14), ack => RPIPE_Block2_start_2065_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2065_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2065_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2065_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2068_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2068_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2068_Sample/rr
      -- 
    ca_5257_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2065_inst_ack_1, ack => convTransposeC_CP_5119_elements(15)); -- 
    rr_5265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(15), ack => RPIPE_Block2_start_2068_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2068_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2068_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2068_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2068_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2068_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2068_Update/cr
      -- 
    ra_5266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2068_inst_ack_0, ack => convTransposeC_CP_5119_elements(16)); -- 
    cr_5270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(16), ack => RPIPE_Block2_start_2068_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2068_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2068_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2068_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2071_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2071_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2071_Sample/rr
      -- 
    ca_5271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2068_inst_ack_1, ack => convTransposeC_CP_5119_elements(17)); -- 
    rr_5279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(17), ack => RPIPE_Block2_start_2071_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2071_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2071_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2071_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2071_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2071_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2071_Update/cr
      -- 
    ra_5280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2071_inst_ack_0, ack => convTransposeC_CP_5119_elements(18)); -- 
    cr_5284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(18), ack => RPIPE_Block2_start_2071_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2071_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2071_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2071_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2074_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2074_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2074_Sample/rr
      -- 
    ca_5285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2071_inst_ack_1, ack => convTransposeC_CP_5119_elements(19)); -- 
    rr_5293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(19), ack => RPIPE_Block2_start_2074_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2074_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2074_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2074_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2074_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2074_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2074_Update/cr
      -- 
    ra_5294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2074_inst_ack_0, ack => convTransposeC_CP_5119_elements(20)); -- 
    cr_5298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(20), ack => RPIPE_Block2_start_2074_inst_req_1); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2074_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2074_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2074_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2077_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2077_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2077_Sample/rr
      -- 
    ca_5299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2074_inst_ack_1, ack => convTransposeC_CP_5119_elements(21)); -- 
    rr_5307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(21), ack => RPIPE_Block2_start_2077_inst_req_0); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2077_Update/cr
      -- CP-element group 22: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2077_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2077_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2077_update_start_
      -- CP-element group 22: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2077_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2077_Sample/ra
      -- 
    ra_5308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2077_inst_ack_0, ack => convTransposeC_CP_5119_elements(22)); -- 
    cr_5312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(22), ack => RPIPE_Block2_start_2077_inst_req_1); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2080_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2077_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2077_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2080_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2080_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2077_update_completed_
      -- 
    ca_5313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2077_inst_ack_1, ack => convTransposeC_CP_5119_elements(23)); -- 
    rr_5321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(23), ack => RPIPE_Block2_start_2080_inst_req_0); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2080_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2080_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2080_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2080_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2080_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2080_Update/cr
      -- 
    ra_5322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2080_inst_ack_0, ack => convTransposeC_CP_5119_elements(24)); -- 
    cr_5326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(24), ack => RPIPE_Block2_start_2080_inst_req_1); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2083_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2080_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2080_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2083_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2083_Sample/rr
      -- CP-element group 25: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2080_Update/$exit
      -- 
    ca_5327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2080_inst_ack_1, ack => convTransposeC_CP_5119_elements(25)); -- 
    rr_5335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(25), ack => RPIPE_Block2_start_2083_inst_req_0); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2083_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2083_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2083_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2083_update_start_
      -- CP-element group 26: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2083_Update/cr
      -- CP-element group 26: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2083_Sample/$exit
      -- 
    ra_5336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2083_inst_ack_0, ack => convTransposeC_CP_5119_elements(26)); -- 
    cr_5340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(26), ack => RPIPE_Block2_start_2083_inst_req_1); -- 
    -- CP-element group 27:  fork  transition  place  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (13) 
      -- CP-element group 27: 	 branch_block_stmt_2045/assign_stmt_2091_to_assign_stmt_2170/type_cast_2100_Update/cr
      -- CP-element group 27: 	 branch_block_stmt_2045/assign_stmt_2091_to_assign_stmt_2170/type_cast_2100_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2083_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2083_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/RPIPE_Block2_start_2083_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_2045/assign_stmt_2091_to_assign_stmt_2170/$entry
      -- CP-element group 27: 	 branch_block_stmt_2045/assign_stmt_2091_to_assign_stmt_2170/type_cast_2100_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_2045/assign_stmt_2091_to_assign_stmt_2170/type_cast_2100_update_start_
      -- CP-element group 27: 	 branch_block_stmt_2045/assign_stmt_2091_to_assign_stmt_2170/type_cast_2100_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_2045/assign_stmt_2091_to_assign_stmt_2170/type_cast_2100_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084__exit__
      -- CP-element group 27: 	 branch_block_stmt_2045/assign_stmt_2091_to_assign_stmt_2170__entry__
      -- CP-element group 27: 	 branch_block_stmt_2045/assign_stmt_2048_to_assign_stmt_2084/$exit
      -- 
    ca_5341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2083_inst_ack_1, ack => convTransposeC_CP_5119_elements(27)); -- 
    cr_5357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(27), ack => type_cast_2100_inst_req_1); -- 
    rr_5352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(27), ack => type_cast_2100_inst_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2045/assign_stmt_2091_to_assign_stmt_2170/type_cast_2100_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2045/assign_stmt_2091_to_assign_stmt_2170/type_cast_2100_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2045/assign_stmt_2091_to_assign_stmt_2170/type_cast_2100_Sample/ra
      -- 
    ra_5353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2100_inst_ack_0, ack => convTransposeC_CP_5119_elements(28)); -- 
    -- CP-element group 29:  fork  transition  place  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	67 
    -- CP-element group 29: 	68 
    -- CP-element group 29: 	70 
    -- CP-element group 29: 	71 
    -- CP-element group 29: 	72 
    -- CP-element group 29:  members (21) 
      -- CP-element group 29: 	 branch_block_stmt_2045/assign_stmt_2091_to_assign_stmt_2170/type_cast_2100_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2045/assign_stmt_2091_to_assign_stmt_2170/type_cast_2100_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_2045/assign_stmt_2091_to_assign_stmt_2170/$exit
      -- CP-element group 29: 	 branch_block_stmt_2045/assign_stmt_2091_to_assign_stmt_2170/type_cast_2100_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2045/assign_stmt_2091_to_assign_stmt_2170__exit__
      -- CP-element group 29: 	 branch_block_stmt_2045/entry_whilex_xbody
      -- CP-element group 29: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 29: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2194/$entry
      -- CP-element group 29: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/$entry
      -- CP-element group 29: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/$entry
      -- CP-element group 29: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/cr
      -- CP-element group 29: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2187/$entry
      -- CP-element group 29: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2180/$entry
      -- CP-element group 29: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2173/$entry
      -- CP-element group 29: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_sources/$entry
      -- 
    ca_5358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2100_inst_ack_1, ack => convTransposeC_CP_5119_elements(29)); -- 
    rr_5748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(29), ack => type_cast_2197_inst_req_0); -- 
    cr_5753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(29), ack => type_cast_2197_inst_req_1); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	92 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2214_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2214_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2214_Sample/ra
      -- 
    ra_5370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2214_inst_ack_0, ack => convTransposeC_CP_5119_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	92 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	44 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2214_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2214_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2214_Update/ca
      -- 
    ca_5375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2214_inst_ack_1, ack => convTransposeC_CP_5119_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	92 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2228_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2228_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2228_sample_completed_
      -- 
    ra_5384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2228_inst_ack_0, ack => convTransposeC_CP_5119_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	92 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	44 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2228_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2228_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2228_Update/ca
      -- 
    ca_5389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2228_inst_ack_1, ack => convTransposeC_CP_5119_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	92 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2242_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2242_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2242_Sample/ra
      -- 
    ra_5398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2242_inst_ack_0, ack => convTransposeC_CP_5119_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	92 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	44 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2242_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2242_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2242_Update/ca
      -- 
    ca_5403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2242_inst_ack_1, ack => convTransposeC_CP_5119_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	92 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2284_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2284_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2284_Sample/ra
      -- 
    ra_5412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2284_inst_ack_0, ack => convTransposeC_CP_5119_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	92 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (16) 
      -- CP-element group 37: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_final_index_sum_regn_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_index_scale_1/scale_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_final_index_sum_regn_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_index_resized_1
      -- CP-element group 37: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_index_scaled_1
      -- CP-element group 37: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_index_computed_1
      -- CP-element group 37: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_index_resize_1/$entry
      -- CP-element group 37: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_index_resize_1/$exit
      -- CP-element group 37: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_index_resize_1/index_resize_req
      -- CP-element group 37: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2284_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_index_resize_1/index_resize_ack
      -- CP-element group 37: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_index_scale_1/$entry
      -- CP-element group 37: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2284_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2284_Update/ca
      -- CP-element group 37: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_index_scale_1/$exit
      -- CP-element group 37: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_index_scale_1/scale_rename_req
      -- 
    ca_5417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2284_inst_ack_1, ack => convTransposeC_CP_5119_elements(37)); -- 
    req_5442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(37), ack => array_obj_ref_2290_index_offset_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	54 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_final_index_sum_regn_sample_complete
      -- CP-element group 38: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_final_index_sum_regn_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_final_index_sum_regn_Sample/$exit
      -- 
    ack_5443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2290_index_offset_ack_0, ack => convTransposeC_CP_5119_elements(38)); -- 
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	92 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (11) 
      -- CP-element group 39: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_final_index_sum_regn_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_final_index_sum_regn_Update/ack
      -- CP-element group 39: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_offset_calculated
      -- CP-element group 39: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2291_request/$entry
      -- CP-element group 39: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2291_request/req
      -- CP-element group 39: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2291_sample_start_
      -- 
    ack_5448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2290_index_offset_ack_1, ack => convTransposeC_CP_5119_elements(39)); -- 
    req_5457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(39), ack => addr_of_2291_final_reg_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2291_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2291_request/$exit
      -- CP-element group 40: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2291_request/ack
      -- 
    ack_5458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2291_final_reg_ack_0, ack => convTransposeC_CP_5119_elements(40)); -- 
    -- CP-element group 41:  join  fork  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	92 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (24) 
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_base_addr_resize/base_resize_req
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Sample/word_access_start/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_base_addr_resize/$exit
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_base_addr_resize/base_resize_ack
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_base_plus_offset/$entry
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2291_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_base_plus_offset/$exit
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_word_addrgen/$entry
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2291_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2291_complete/ack
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_word_addrgen/$exit
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Sample/word_access_start/word_0/rr
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_word_addrgen/root_register_req
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_base_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_word_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_base_address_resized
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_word_addrgen/root_register_ack
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Sample/word_access_start/$entry
      -- CP-element group 41: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_base_addr_resize/$entry
      -- 
    ack_5463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2291_final_reg_ack_1, ack => convTransposeC_CP_5119_elements(41)); -- 
    rr_5496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(41), ack => ptr_deref_2295_load_0_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Sample/word_access_start/$exit
      -- CP-element group 42: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Sample/word_access_start/word_0/$exit
      -- CP-element group 42: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Sample/word_access_start/word_0/ra
      -- CP-element group 42: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Sample/$exit
      -- 
    ra_5497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_load_0_ack_0, ack => convTransposeC_CP_5119_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	92 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	51 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Update/word_access_complete/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Update/word_access_complete/word_0/ca
      -- CP-element group 43: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Update/ptr_deref_2295_Merge/$entry
      -- CP-element group 43: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Update/ptr_deref_2295_Merge/$exit
      -- CP-element group 43: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Update/ptr_deref_2295_Merge/merge_req
      -- CP-element group 43: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Update/ptr_deref_2295_Merge/merge_ack
      -- CP-element group 43: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Update/word_access_complete/$exit
      -- 
    ca_5508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2295_load_0_ack_1, ack => convTransposeC_CP_5119_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	31 
    -- CP-element group 44: 	33 
    -- CP-element group 44: 	35 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2305_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2305_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2305_Sample/rr
      -- 
    rr_5521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(44), ack => type_cast_2305_inst_req_0); -- 
    convTransposeC_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(31) & convTransposeC_CP_5119_elements(33) & convTransposeC_CP_5119_elements(35);
      gj_convTransposeC_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2305_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2305_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2305_Sample/ra
      -- 
    ra_5522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2305_inst_ack_0, ack => convTransposeC_CP_5119_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	92 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (16) 
      -- CP-element group 46: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_final_index_sum_regn_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2305_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2305_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2305_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_index_resized_1
      -- CP-element group 46: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_final_index_sum_regn_Sample/req
      -- CP-element group 46: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_index_scaled_1
      -- CP-element group 46: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_index_computed_1
      -- CP-element group 46: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_index_resize_1/$entry
      -- CP-element group 46: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_index_resize_1/$exit
      -- CP-element group 46: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_index_resize_1/index_resize_req
      -- CP-element group 46: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_index_resize_1/index_resize_ack
      -- CP-element group 46: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_index_scale_1/$entry
      -- CP-element group 46: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_index_scale_1/$exit
      -- CP-element group 46: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_index_scale_1/scale_rename_req
      -- CP-element group 46: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_index_scale_1/scale_rename_ack
      -- 
    ca_5527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2305_inst_ack_1, ack => convTransposeC_CP_5119_elements(46)); -- 
    req_5552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(46), ack => array_obj_ref_2311_index_offset_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	54 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_final_index_sum_regn_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_final_index_sum_regn_sample_complete
      -- CP-element group 47: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_final_index_sum_regn_Sample/ack
      -- 
    ack_5553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2311_index_offset_ack_0, ack => convTransposeC_CP_5119_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	92 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (11) 
      -- CP-element group 48: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_root_address_calculated
      -- CP-element group 48: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_final_index_sum_regn_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2312_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_offset_calculated
      -- CP-element group 48: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2312_request/$entry
      -- CP-element group 48: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_base_plus_offset/sum_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2312_request/req
      -- CP-element group 48: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_base_plus_offset/sum_rename_req
      -- CP-element group 48: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_base_plus_offset/$entry
      -- CP-element group 48: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_base_plus_offset/$exit
      -- CP-element group 48: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_final_index_sum_regn_Update/ack
      -- 
    ack_5558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2311_index_offset_ack_1, ack => convTransposeC_CP_5119_elements(48)); -- 
    req_5567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(48), ack => addr_of_2312_final_reg_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2312_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2312_request/$exit
      -- CP-element group 49: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2312_request/ack
      -- 
    ack_5568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2312_final_reg_ack_0, ack => convTransposeC_CP_5119_elements(49)); -- 
    -- CP-element group 50:  fork  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	92 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (19) 
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_word_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2312_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_base_address_resized
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_base_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2312_complete/ack
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_base_addr_resize/$entry
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_base_addr_resize/$exit
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_base_addr_resize/base_resize_req
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_base_addr_resize/base_resize_ack
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_base_plus_offset/sum_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2312_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_word_addrgen/$entry
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_word_addrgen/$exit
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_word_addrgen/root_register_req
      -- CP-element group 50: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_word_addrgen/root_register_ack
      -- 
    ack_5573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2312_final_reg_ack_1, ack => convTransposeC_CP_5119_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	43 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Sample/ptr_deref_2315_Split/$entry
      -- CP-element group 51: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Sample/ptr_deref_2315_Split/$exit
      -- CP-element group 51: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Sample/ptr_deref_2315_Split/split_req
      -- CP-element group 51: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Sample/ptr_deref_2315_Split/split_ack
      -- CP-element group 51: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Sample/word_access_start/word_0/rr
      -- 
    rr_5611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(51), ack => ptr_deref_2315_store_0_req_0); -- 
    convTransposeC_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(43) & convTransposeC_CP_5119_elements(50);
      gj_convTransposeC_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Sample/word_access_start/word_0/ra
      -- 
    ra_5612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2315_store_0_ack_0, ack => convTransposeC_CP_5119_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	92 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Update/word_access_complete/word_0/ca
      -- 
    ca_5623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2315_store_0_ack_1, ack => convTransposeC_CP_5119_elements(53)); -- 
    -- CP-element group 54:  branch  join  transition  place  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	38 
    -- CP-element group 54: 	47 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (10) 
      -- CP-element group 54: 	 branch_block_stmt_2045/R_cmp_2330_place
      -- CP-element group 54: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/$exit
      -- CP-element group 54: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328__exit__
      -- CP-element group 54: 	 branch_block_stmt_2045/if_stmt_2329__entry__
      -- CP-element group 54: 	 branch_block_stmt_2045/if_stmt_2329_dead_link/$entry
      -- CP-element group 54: 	 branch_block_stmt_2045/if_stmt_2329_eval_test/$entry
      -- CP-element group 54: 	 branch_block_stmt_2045/if_stmt_2329_eval_test/$exit
      -- CP-element group 54: 	 branch_block_stmt_2045/if_stmt_2329_eval_test/branch_req
      -- CP-element group 54: 	 branch_block_stmt_2045/if_stmt_2329_if_link/$entry
      -- CP-element group 54: 	 branch_block_stmt_2045/if_stmt_2329_else_link/$entry
      -- 
    branch_req_5631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(54), ack => if_stmt_2329_branch_req_0); -- 
    convTransposeC_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(38) & convTransposeC_CP_5119_elements(47) & convTransposeC_CP_5119_elements(53);
      gj_convTransposeC_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	101 
    -- CP-element group 55: 	102 
    -- CP-element group 55: 	104 
    -- CP-element group 55: 	105 
    -- CP-element group 55: 	107 
    -- CP-element group 55: 	108 
    -- CP-element group 55:  members (40) 
      -- CP-element group 55: 	 branch_block_stmt_2045/whilex_xbody_ifx_xthen
      -- CP-element group 55: 	 branch_block_stmt_2045/merge_stmt_2335__exit__
      -- CP-element group 55: 	 branch_block_stmt_2045/assign_stmt_2341__entry__
      -- CP-element group 55: 	 branch_block_stmt_2045/assign_stmt_2341__exit__
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139
      -- CP-element group 55: 	 branch_block_stmt_2045/if_stmt_2329_if_link/$exit
      -- CP-element group 55: 	 branch_block_stmt_2045/if_stmt_2329_if_link/if_choice_transition
      -- CP-element group 55: 	 branch_block_stmt_2045/assign_stmt_2341/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/assign_stmt_2341/$exit
      -- CP-element group 55: 	 branch_block_stmt_2045/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 55: 	 branch_block_stmt_2045/merge_stmt_2335_PhiReqMerge
      -- CP-element group 55: 	 branch_block_stmt_2045/merge_stmt_2335_PhiAck/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/merge_stmt_2335_PhiAck/$exit
      -- CP-element group 55: 	 branch_block_stmt_2045/merge_stmt_2335_PhiAck/dummy
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2391/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_sources/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_sources/type_cast_2397/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_sources/type_cast_2397/SplitProtocol/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_sources/type_cast_2397/SplitProtocol/Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_sources/type_cast_2397/SplitProtocol/Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_sources/type_cast_2397/SplitProtocol/Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_sources/type_cast_2397/SplitProtocol/Update/cr
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2398/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2403/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2403/SplitProtocol/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2403/SplitProtocol/Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2403/SplitProtocol/Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2403/SplitProtocol/Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2403/SplitProtocol/Update/cr
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2404/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2409/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2409/SplitProtocol/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2409/SplitProtocol/Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2409/SplitProtocol/Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2409/SplitProtocol/Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2409/SplitProtocol/Update/cr
      -- 
    if_choice_transition_5636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2329_branch_ack_1, ack => convTransposeC_CP_5119_elements(55)); -- 
    rr_5982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(55), ack => type_cast_2397_inst_req_0); -- 
    cr_5987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(55), ack => type_cast_2397_inst_req_1); -- 
    rr_6005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(55), ack => type_cast_2403_inst_req_0); -- 
    cr_6010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(55), ack => type_cast_2403_inst_req_1); -- 
    rr_6028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(55), ack => type_cast_2409_inst_req_0); -- 
    cr_6033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(55), ack => type_cast_2409_inst_req_1); -- 
    -- CP-element group 56:  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	58 
    -- CP-element group 56: 	60 
    -- CP-element group 56: 	62 
    -- CP-element group 56:  members (24) 
      -- CP-element group 56: 	 branch_block_stmt_2045/whilex_xbody_ifx_xelse
      -- CP-element group 56: 	 branch_block_stmt_2045/merge_stmt_2343__exit__
      -- CP-element group 56: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383__entry__
      -- CP-element group 56: 	 branch_block_stmt_2045/if_stmt_2329_else_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_2045/if_stmt_2329_else_link/else_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/$entry
      -- CP-element group 56: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2352_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2352_update_start_
      -- CP-element group 56: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2352_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2352_Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2352_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2352_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2361_update_start_
      -- CP-element group 56: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2361_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2361_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2377_update_start_
      -- CP-element group 56: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2377_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2377_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_2045/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_2045/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_2045/merge_stmt_2343_PhiReqMerge
      -- CP-element group 56: 	 branch_block_stmt_2045/merge_stmt_2343_PhiAck/$entry
      -- CP-element group 56: 	 branch_block_stmt_2045/merge_stmt_2343_PhiAck/$exit
      -- CP-element group 56: 	 branch_block_stmt_2045/merge_stmt_2343_PhiAck/dummy
      -- 
    else_choice_transition_5640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2329_branch_ack_0, ack => convTransposeC_CP_5119_elements(56)); -- 
    rr_5656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(56), ack => type_cast_2352_inst_req_0); -- 
    cr_5661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(56), ack => type_cast_2352_inst_req_1); -- 
    cr_5675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(56), ack => type_cast_2361_inst_req_1); -- 
    cr_5689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(56), ack => type_cast_2377_inst_req_1); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2352_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2352_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2352_Sample/ra
      -- 
    ra_5657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2352_inst_ack_0, ack => convTransposeC_CP_5119_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2352_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2352_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2352_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2361_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2361_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2361_Sample/rr
      -- 
    ca_5662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2352_inst_ack_1, ack => convTransposeC_CP_5119_elements(58)); -- 
    rr_5670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(58), ack => type_cast_2361_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2361_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2361_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2361_Sample/ra
      -- 
    ra_5671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2361_inst_ack_0, ack => convTransposeC_CP_5119_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	56 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2361_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2361_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2361_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2377_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2377_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2377_Sample/rr
      -- 
    ca_5676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2361_inst_ack_1, ack => convTransposeC_CP_5119_elements(60)); -- 
    rr_5684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(60), ack => type_cast_2377_inst_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2377_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2377_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2377_Sample/ra
      -- 
    ra_5685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2377_inst_ack_0, ack => convTransposeC_CP_5119_elements(61)); -- 
    -- CP-element group 62:  branch  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	56 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (13) 
      -- CP-element group 62: 	 branch_block_stmt_2045/R_cmp128_2385_place
      -- CP-element group 62: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383__exit__
      -- CP-element group 62: 	 branch_block_stmt_2045/if_stmt_2384__entry__
      -- CP-element group 62: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/$exit
      -- CP-element group 62: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2377_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2377_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_2045/assign_stmt_2349_to_assign_stmt_2383/type_cast_2377_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_2045/if_stmt_2384_dead_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_2045/if_stmt_2384_eval_test/$entry
      -- CP-element group 62: 	 branch_block_stmt_2045/if_stmt_2384_eval_test/$exit
      -- CP-element group 62: 	 branch_block_stmt_2045/if_stmt_2384_eval_test/branch_req
      -- CP-element group 62: 	 branch_block_stmt_2045/if_stmt_2384_if_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_2045/if_stmt_2384_else_link/$entry
      -- 
    ca_5690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2377_inst_ack_1, ack => convTransposeC_CP_5119_elements(62)); -- 
    branch_req_5698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(62), ack => if_stmt_2384_branch_req_0); -- 
    -- CP-element group 63:  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (15) 
      -- CP-element group 63: 	 branch_block_stmt_2045/ifx_xelse_whilex_xend
      -- CP-element group 63: 	 branch_block_stmt_2045/merge_stmt_2418__exit__
      -- CP-element group 63: 	 branch_block_stmt_2045/assign_stmt_2423__entry__
      -- CP-element group 63: 	 branch_block_stmt_2045/if_stmt_2384_if_link/$exit
      -- CP-element group 63: 	 branch_block_stmt_2045/if_stmt_2384_if_link/if_choice_transition
      -- CP-element group 63: 	 branch_block_stmt_2045/assign_stmt_2423/$entry
      -- CP-element group 63: 	 branch_block_stmt_2045/assign_stmt_2423/WPIPE_Block2_done_2420_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_2045/assign_stmt_2423/WPIPE_Block2_done_2420_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_2045/assign_stmt_2423/WPIPE_Block2_done_2420_Sample/req
      -- CP-element group 63: 	 branch_block_stmt_2045/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 63: 	 branch_block_stmt_2045/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 63: 	 branch_block_stmt_2045/merge_stmt_2418_PhiReqMerge
      -- CP-element group 63: 	 branch_block_stmt_2045/merge_stmt_2418_PhiAck/$entry
      -- CP-element group 63: 	 branch_block_stmt_2045/merge_stmt_2418_PhiAck/$exit
      -- CP-element group 63: 	 branch_block_stmt_2045/merge_stmt_2418_PhiAck/dummy
      -- 
    if_choice_transition_5703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2384_branch_ack_1, ack => convTransposeC_CP_5119_elements(63)); -- 
    req_5723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(63), ack => WPIPE_Block2_done_2420_inst_req_0); -- 
    -- CP-element group 64:  fork  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	93 
    -- CP-element group 64: 	94 
    -- CP-element group 64: 	95 
    -- CP-element group 64: 	97 
    -- CP-element group 64: 	98 
    -- CP-element group 64:  members (22) 
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139
      -- CP-element group 64: 	 branch_block_stmt_2045/if_stmt_2384_else_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_2045/if_stmt_2384_else_link/else_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2391/$entry
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_sources/$entry
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2398/$entry
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/$entry
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2401/$entry
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2401/SplitProtocol/$entry
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2401/SplitProtocol/Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2401/SplitProtocol/Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2401/SplitProtocol/Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2401/SplitProtocol/Update/cr
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2404/$entry
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/$entry
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2407/$entry
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2407/SplitProtocol/$entry
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2407/SplitProtocol/Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2407/SplitProtocol/Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2407/SplitProtocol/Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2407/SplitProtocol/Update/cr
      -- 
    else_choice_transition_5707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2384_branch_ack_0, ack => convTransposeC_CP_5119_elements(64)); -- 
    rr_5933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(64), ack => type_cast_2401_inst_req_0); -- 
    cr_5938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(64), ack => type_cast_2401_inst_req_1); -- 
    rr_5956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(64), ack => type_cast_2407_inst_req_0); -- 
    cr_5961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(64), ack => type_cast_2407_inst_req_1); -- 
    -- CP-element group 65:  transition  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (6) 
      -- CP-element group 65: 	 branch_block_stmt_2045/assign_stmt_2423/WPIPE_Block2_done_2420_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_2045/assign_stmt_2423/WPIPE_Block2_done_2420_update_start_
      -- CP-element group 65: 	 branch_block_stmt_2045/assign_stmt_2423/WPIPE_Block2_done_2420_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_2045/assign_stmt_2423/WPIPE_Block2_done_2420_Sample/ack
      -- CP-element group 65: 	 branch_block_stmt_2045/assign_stmt_2423/WPIPE_Block2_done_2420_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_2045/assign_stmt_2423/WPIPE_Block2_done_2420_Update/req
      -- 
    ack_5724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2420_inst_ack_0, ack => convTransposeC_CP_5119_elements(65)); -- 
    req_5728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(65), ack => WPIPE_Block2_done_2420_inst_req_1); -- 
    -- CP-element group 66:  transition  place  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (16) 
      -- CP-element group 66: 	 $exit
      -- CP-element group 66: 	 branch_block_stmt_2045/$exit
      -- CP-element group 66: 	 branch_block_stmt_2045/branch_block_stmt_2045__exit__
      -- CP-element group 66: 	 branch_block_stmt_2045/assign_stmt_2423__exit__
      -- CP-element group 66: 	 branch_block_stmt_2045/return__
      -- CP-element group 66: 	 branch_block_stmt_2045/merge_stmt_2425__exit__
      -- CP-element group 66: 	 branch_block_stmt_2045/assign_stmt_2423/$exit
      -- CP-element group 66: 	 branch_block_stmt_2045/assign_stmt_2423/WPIPE_Block2_done_2420_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_2045/assign_stmt_2423/WPIPE_Block2_done_2420_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_2045/assign_stmt_2423/WPIPE_Block2_done_2420_Update/ack
      -- CP-element group 66: 	 branch_block_stmt_2045/return___PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_2045/return___PhiReq/$exit
      -- CP-element group 66: 	 branch_block_stmt_2045/merge_stmt_2425_PhiReqMerge
      -- CP-element group 66: 	 branch_block_stmt_2045/merge_stmt_2425_PhiAck/$entry
      -- CP-element group 66: 	 branch_block_stmt_2045/merge_stmt_2425_PhiAck/$exit
      -- CP-element group 66: 	 branch_block_stmt_2045/merge_stmt_2425_PhiAck/dummy
      -- 
    ack_5729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2420_inst_ack_1, ack => convTransposeC_CP_5119_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	29 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Sample/ra
      -- 
    ra_5749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2197_inst_ack_0, ack => convTransposeC_CP_5119_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	29 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/Update/ca
      -- 
    ca_5754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2197_inst_ack_1, ack => convTransposeC_CP_5119_elements(68)); -- 
    -- CP-element group 69:  join  transition  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	73 
    -- CP-element group 69:  members (5) 
      -- CP-element group 69: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2194/$exit
      -- CP-element group 69: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/$exit
      -- CP-element group 69: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/$exit
      -- CP-element group 69: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2197/SplitProtocol/$exit
      -- CP-element group 69: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_req
      -- 
    phi_stmt_2194_req_5755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2194_req_5755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(69), ack => phi_stmt_2194_req_0); -- 
    convTransposeC_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(67) & convTransposeC_CP_5119_elements(68);
      gj_convTransposeC_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  output  delay-element  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	29 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	73 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2187/$exit
      -- CP-element group 70: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/$exit
      -- CP-element group 70: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2193_konst_delay_trans
      -- CP-element group 70: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_req
      -- 
    phi_stmt_2187_req_5763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2187_req_5763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(70), ack => phi_stmt_2187_req_1); -- 
    -- Element group convTransposeC_CP_5119_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => convTransposeC_CP_5119_elements(29), ack => convTransposeC_CP_5119_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  transition  output  delay-element  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	29 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2180/$exit
      -- CP-element group 71: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_sources/$exit
      -- CP-element group 71: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_sources/type_cast_2184_konst_delay_trans
      -- CP-element group 71: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_req
      -- 
    phi_stmt_2180_req_5771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2180_req_5771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(71), ack => phi_stmt_2180_req_0); -- 
    -- Element group convTransposeC_CP_5119_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => convTransposeC_CP_5119_elements(29), ack => convTransposeC_CP_5119_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  transition  output  delay-element  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	29 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2173/$exit
      -- CP-element group 72: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_sources/$exit
      -- CP-element group 72: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_sources/type_cast_2177_konst_delay_trans
      -- CP-element group 72: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_req
      -- 
    phi_stmt_2173_req_5779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2173_req_5779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(72), ack => phi_stmt_2173_req_0); -- 
    -- Element group convTransposeC_CP_5119_elements(72) is a control-delay.
    cp_element_72_delay: control_delay_element  generic map(name => " 72_delay", delay_value => 1)  port map(req => convTransposeC_CP_5119_elements(29), ack => convTransposeC_CP_5119_elements(72), clk => clk, reset =>reset);
    -- CP-element group 73:  join  transition  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	69 
    -- CP-element group 73: 	70 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	87 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_2045/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(69) & convTransposeC_CP_5119_elements(70) & convTransposeC_CP_5119_elements(71) & convTransposeC_CP_5119_elements(72);
      gj_convTransposeC_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	1 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Sample/ra
      -- 
    ra_5799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2199_inst_ack_0, ack => convTransposeC_CP_5119_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	1 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/Update/ca
      -- 
    ca_5804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2199_inst_ack_1, ack => convTransposeC_CP_5119_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	86 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2194/$exit
      -- CP-element group 76: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/$exit
      -- CP-element group 76: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_sources/type_cast_2199/SplitProtocol/$exit
      -- CP-element group 76: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2194/phi_stmt_2194_req
      -- 
    phi_stmt_2194_req_5805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2194_req_5805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(76), ack => phi_stmt_2194_req_1); -- 
    convTransposeC_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(74) & convTransposeC_CP_5119_elements(75);
      gj_convTransposeC_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	1 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2190/SplitProtocol/Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2190/SplitProtocol/Sample/ra
      -- 
    ra_5822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2190_inst_ack_0, ack => convTransposeC_CP_5119_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	1 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2190/SplitProtocol/Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2190/SplitProtocol/Update/ca
      -- 
    ca_5827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2190_inst_ack_1, ack => convTransposeC_CP_5119_elements(78)); -- 
    -- CP-element group 79:  join  transition  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	86 
    -- CP-element group 79:  members (5) 
      -- CP-element group 79: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2187/$exit
      -- CP-element group 79: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2190/$exit
      -- CP-element group 79: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_sources/type_cast_2190/SplitProtocol/$exit
      -- CP-element group 79: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2187/phi_stmt_2187_req
      -- 
    phi_stmt_2187_req_5828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2187_req_5828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(79), ack => phi_stmt_2187_req_0); -- 
    convTransposeC_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(77) & convTransposeC_CP_5119_elements(78);
      gj_convTransposeC_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	1 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_sources/type_cast_2186/SplitProtocol/Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_sources/type_cast_2186/SplitProtocol/Sample/ra
      -- 
    ra_5845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2186_inst_ack_0, ack => convTransposeC_CP_5119_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	1 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_sources/type_cast_2186/SplitProtocol/Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_sources/type_cast_2186/SplitProtocol/Update/ca
      -- 
    ca_5850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2186_inst_ack_1, ack => convTransposeC_CP_5119_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	86 
    -- CP-element group 82:  members (5) 
      -- CP-element group 82: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2180/$exit
      -- CP-element group 82: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_sources/type_cast_2186/$exit
      -- CP-element group 82: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_sources/type_cast_2186/SplitProtocol/$exit
      -- CP-element group 82: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2180/phi_stmt_2180_req
      -- 
    phi_stmt_2180_req_5851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2180_req_5851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(82), ack => phi_stmt_2180_req_1); -- 
    convTransposeC_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(80) & convTransposeC_CP_5119_elements(81);
      gj_convTransposeC_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	1 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_sources/type_cast_2179/SplitProtocol/Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_sources/type_cast_2179/SplitProtocol/Sample/ra
      -- 
    ra_5868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2179_inst_ack_0, ack => convTransposeC_CP_5119_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	1 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_sources/type_cast_2179/SplitProtocol/Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_sources/type_cast_2179/SplitProtocol/Update/ca
      -- 
    ca_5873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2179_inst_ack_1, ack => convTransposeC_CP_5119_elements(84)); -- 
    -- CP-element group 85:  join  transition  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2173/$exit
      -- CP-element group 85: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_sources/$exit
      -- CP-element group 85: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_sources/type_cast_2179/$exit
      -- CP-element group 85: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_sources/type_cast_2179/SplitProtocol/$exit
      -- CP-element group 85: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/phi_stmt_2173/phi_stmt_2173_req
      -- 
    phi_stmt_2173_req_5874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2173_req_5874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(85), ack => phi_stmt_2173_req_1); -- 
    convTransposeC_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(83) & convTransposeC_CP_5119_elements(84);
      gj_convTransposeC_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  join  transition  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	76 
    -- CP-element group 86: 	79 
    -- CP-element group 86: 	82 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_2045/ifx_xend139_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(76) & convTransposeC_CP_5119_elements(79) & convTransposeC_CP_5119_elements(82) & convTransposeC_CP_5119_elements(85);
      gj_convTransposeC_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  merge  fork  transition  place  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	73 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	89 
    -- CP-element group 87: 	90 
    -- CP-element group 87: 	91 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2045/merge_stmt_2172_PhiReqMerge
      -- CP-element group 87: 	 branch_block_stmt_2045/merge_stmt_2172_PhiAck/$entry
      -- 
    convTransposeC_CP_5119_elements(87) <= OrReduce(convTransposeC_CP_5119_elements(73) & convTransposeC_CP_5119_elements(86));
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	92 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_2045/merge_stmt_2172_PhiAck/phi_stmt_2173_ack
      -- 
    phi_stmt_2173_ack_5879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2173_ack_0, ack => convTransposeC_CP_5119_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	92 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_2045/merge_stmt_2172_PhiAck/phi_stmt_2180_ack
      -- 
    phi_stmt_2180_ack_5880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2180_ack_0, ack => convTransposeC_CP_5119_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_2045/merge_stmt_2172_PhiAck/phi_stmt_2187_ack
      -- 
    phi_stmt_2187_ack_5881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2187_ack_0, ack => convTransposeC_CP_5119_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	87 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_2045/merge_stmt_2172_PhiAck/phi_stmt_2194_ack
      -- 
    phi_stmt_2194_ack_5882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2194_ack_0, ack => convTransposeC_CP_5119_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  place  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	88 
    -- CP-element group 92: 	89 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	30 
    -- CP-element group 92: 	31 
    -- CP-element group 92: 	32 
    -- CP-element group 92: 	33 
    -- CP-element group 92: 	34 
    -- CP-element group 92: 	35 
    -- CP-element group 92: 	36 
    -- CP-element group 92: 	37 
    -- CP-element group 92: 	39 
    -- CP-element group 92: 	41 
    -- CP-element group 92: 	43 
    -- CP-element group 92: 	46 
    -- CP-element group 92: 	48 
    -- CP-element group 92: 	50 
    -- CP-element group 92: 	53 
    -- CP-element group 92:  members (53) 
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2228_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_final_index_sum_regn_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_final_index_sum_regn_Update/req
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2290_final_index_sum_regn_update_start
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2291_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2228_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2228_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Update/word_access_complete/word_0/cr
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2228_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2214_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2228_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2305_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2242_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2214_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2305_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2305_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2242_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2291_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2312_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2291_complete/req
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2242_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2242_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2242_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2214_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2214_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2242_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2284_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2284_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2214_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2284_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2284_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2214_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2284_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2312_complete/req
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2228_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/type_cast_2284_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_final_index_sum_regn_update_start
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_final_index_sum_regn_Update/req
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Update/word_access_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/array_obj_ref_2311_final_index_sum_regn_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/addr_of_2312_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/merge_stmt_2172__exit__
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328__entry__
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2295_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Update/word_access_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_2045/assign_stmt_2206_to_assign_stmt_2328/ptr_deref_2315_Update/word_access_complete/word_0/cr
      -- CP-element group 92: 	 branch_block_stmt_2045/merge_stmt_2172_PhiAck/$exit
      -- 
    req_5447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(92), ack => array_obj_ref_2290_index_offset_req_1); -- 
    rr_5383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(92), ack => type_cast_2228_inst_req_0); -- 
    cr_5507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(92), ack => ptr_deref_2295_load_0_req_1); -- 
    cr_5388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(92), ack => type_cast_2228_inst_req_1); -- 
    cr_5526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(92), ack => type_cast_2305_inst_req_1); -- 
    req_5462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(92), ack => addr_of_2291_final_reg_req_1); -- 
    rr_5397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(92), ack => type_cast_2242_inst_req_0); -- 
    rr_5369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(92), ack => type_cast_2214_inst_req_0); -- 
    cr_5402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(92), ack => type_cast_2242_inst_req_1); -- 
    rr_5411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(92), ack => type_cast_2284_inst_req_0); -- 
    cr_5374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(92), ack => type_cast_2214_inst_req_1); -- 
    req_5572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(92), ack => addr_of_2312_final_reg_req_1); -- 
    cr_5416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(92), ack => type_cast_2284_inst_req_1); -- 
    req_5557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(92), ack => array_obj_ref_2311_index_offset_req_1); -- 
    cr_5622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(92), ack => ptr_deref_2315_store_0_req_1); -- 
    convTransposeC_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(88) & convTransposeC_CP_5119_elements(89) & convTransposeC_CP_5119_elements(90) & convTransposeC_CP_5119_elements(91);
      gj_convTransposeC_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  output  delay-element  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	64 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	100 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2391/$exit
      -- CP-element group 93: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_sources/type_cast_2395_konst_delay_trans
      -- CP-element group 93: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_req
      -- 
    phi_stmt_2391_req_5917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2391_req_5917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(93), ack => phi_stmt_2391_req_0); -- 
    -- Element group convTransposeC_CP_5119_elements(93) is a control-delay.
    cp_element_93_delay: control_delay_element  generic map(name => " 93_delay", delay_value => 1)  port map(req => convTransposeC_CP_5119_elements(64), ack => convTransposeC_CP_5119_elements(93), clk => clk, reset =>reset);
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	64 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2401/SplitProtocol/Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2401/SplitProtocol/Sample/ra
      -- 
    ra_5934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2401_inst_ack_0, ack => convTransposeC_CP_5119_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	64 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2401/SplitProtocol/Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2401/SplitProtocol/Update/ca
      -- 
    ca_5939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2401_inst_ack_1, ack => convTransposeC_CP_5119_elements(95)); -- 
    -- CP-element group 96:  join  transition  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	100 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2398/$exit
      -- CP-element group 96: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/$exit
      -- CP-element group 96: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2401/$exit
      -- CP-element group 96: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2401/SplitProtocol/$exit
      -- CP-element group 96: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_req
      -- 
    phi_stmt_2398_req_5940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2398_req_5940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(96), ack => phi_stmt_2398_req_0); -- 
    convTransposeC_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(94) & convTransposeC_CP_5119_elements(95);
      gj_convTransposeC_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	64 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2407/SplitProtocol/Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2407/SplitProtocol/Sample/ra
      -- 
    ra_5957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2407_inst_ack_0, ack => convTransposeC_CP_5119_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	64 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2407/SplitProtocol/Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2407/SplitProtocol/Update/ca
      -- 
    ca_5962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2407_inst_ack_1, ack => convTransposeC_CP_5119_elements(98)); -- 
    -- CP-element group 99:  join  transition  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2404/$exit
      -- CP-element group 99: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/$exit
      -- CP-element group 99: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2407/$exit
      -- CP-element group 99: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2407/SplitProtocol/$exit
      -- CP-element group 99: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_req
      -- 
    phi_stmt_2404_req_5963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2404_req_5963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(99), ack => phi_stmt_2404_req_0); -- 
    convTransposeC_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(97) & convTransposeC_CP_5119_elements(98);
      gj_convTransposeC_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  join  transition  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	93 
    -- CP-element group 100: 	96 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	111 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_2045/ifx_xelse_ifx_xend139_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(93) & convTransposeC_CP_5119_elements(96) & convTransposeC_CP_5119_elements(99);
      gj_convTransposeC_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	55 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_sources/type_cast_2397/SplitProtocol/Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_sources/type_cast_2397/SplitProtocol/Sample/ra
      -- 
    ra_5983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2397_inst_ack_0, ack => convTransposeC_CP_5119_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	55 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_sources/type_cast_2397/SplitProtocol/Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_sources/type_cast_2397/SplitProtocol/Update/ca
      -- 
    ca_5988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2397_inst_ack_1, ack => convTransposeC_CP_5119_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	110 
    -- CP-element group 103:  members (5) 
      -- CP-element group 103: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2391/$exit
      -- CP-element group 103: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_sources/$exit
      -- CP-element group 103: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_sources/type_cast_2397/$exit
      -- CP-element group 103: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_sources/type_cast_2397/SplitProtocol/$exit
      -- CP-element group 103: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2391/phi_stmt_2391_req
      -- 
    phi_stmt_2391_req_5989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2391_req_5989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(103), ack => phi_stmt_2391_req_1); -- 
    convTransposeC_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(101) & convTransposeC_CP_5119_elements(102);
      gj_convTransposeC_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	55 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2403/SplitProtocol/Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2403/SplitProtocol/Sample/ra
      -- 
    ra_6006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2403_inst_ack_0, ack => convTransposeC_CP_5119_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	55 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2403/SplitProtocol/Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2403/SplitProtocol/Update/ca
      -- 
    ca_6011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2403_inst_ack_1, ack => convTransposeC_CP_5119_elements(105)); -- 
    -- CP-element group 106:  join  transition  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	110 
    -- CP-element group 106:  members (5) 
      -- CP-element group 106: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2398/$exit
      -- CP-element group 106: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/$exit
      -- CP-element group 106: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2403/$exit
      -- CP-element group 106: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_sources/type_cast_2403/SplitProtocol/$exit
      -- CP-element group 106: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2398/phi_stmt_2398_req
      -- 
    phi_stmt_2398_req_6012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2398_req_6012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(106), ack => phi_stmt_2398_req_1); -- 
    convTransposeC_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(104) & convTransposeC_CP_5119_elements(105);
      gj_convTransposeC_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	55 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2409/SplitProtocol/Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2409/SplitProtocol/Sample/ra
      -- 
    ra_6029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2409_inst_ack_0, ack => convTransposeC_CP_5119_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	55 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2409/SplitProtocol/Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2409/SplitProtocol/Update/ca
      -- 
    ca_6034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2409_inst_ack_1, ack => convTransposeC_CP_5119_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2404/$exit
      -- CP-element group 109: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/$exit
      -- CP-element group 109: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2409/$exit
      -- CP-element group 109: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_sources/type_cast_2409/SplitProtocol/$exit
      -- CP-element group 109: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/phi_stmt_2404/phi_stmt_2404_req
      -- 
    phi_stmt_2404_req_6035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2404_req_6035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_5119_elements(109), ack => phi_stmt_2404_req_1); -- 
    convTransposeC_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(107) & convTransposeC_CP_5119_elements(108);
      gj_convTransposeC_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  transition  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	103 
    -- CP-element group 110: 	106 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_2045/ifx_xthen_ifx_xend139_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(103) & convTransposeC_CP_5119_elements(106) & convTransposeC_CP_5119_elements(109);
      gj_convTransposeC_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  merge  fork  transition  place  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	100 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	113 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_2045/merge_stmt_2390_PhiReqMerge
      -- CP-element group 111: 	 branch_block_stmt_2045/merge_stmt_2390_PhiAck/$entry
      -- 
    convTransposeC_CP_5119_elements(111) <= OrReduce(convTransposeC_CP_5119_elements(100) & convTransposeC_CP_5119_elements(110));
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	115 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2045/merge_stmt_2390_PhiAck/phi_stmt_2391_ack
      -- 
    phi_stmt_2391_ack_6040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2391_ack_0, ack => convTransposeC_CP_5119_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_2045/merge_stmt_2390_PhiAck/phi_stmt_2398_ack
      -- 
    phi_stmt_2398_ack_6041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2398_ack_0, ack => convTransposeC_CP_5119_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_2045/merge_stmt_2390_PhiAck/phi_stmt_2404_ack
      -- 
    phi_stmt_2404_ack_6042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2404_ack_0, ack => convTransposeC_CP_5119_elements(114)); -- 
    -- CP-element group 115:  join  transition  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	112 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	1 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_2045/merge_stmt_2390_PhiAck/$exit
      -- 
    convTransposeC_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeC_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeC_CP_5119_elements(112) & convTransposeC_CP_5119_elements(113) & convTransposeC_CP_5119_elements(114);
      gj_convTransposeC_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_5119_elements(115), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom92_2310_resized : std_logic_vector(13 downto 0);
    signal R_idxprom92_2310_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2289_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2289_scaled : std_logic_vector(13 downto 0);
    signal add104_2341 : std_logic_vector(15 downto 0);
    signal add127_2170 : std_logic_vector(31 downto 0);
    signal add64_2124 : std_logic_vector(31 downto 0);
    signal add83_2265 : std_logic_vector(31 downto 0);
    signal add85_2275 : std_logic_vector(31 downto 0);
    signal add97_2323 : std_logic_vector(31 downto 0);
    signal add_2113 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2211 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2290_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2290_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2290_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2290_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2290_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2290_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2311_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2311_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2311_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2311_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2311_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2311_root_address : std_logic_vector(13 downto 0);
    signal arrayidx88_2292 : std_logic_vector(31 downto 0);
    signal arrayidx93_2313 : std_logic_vector(31 downto 0);
    signal call10_2060 : std_logic_vector(31 downto 0);
    signal call13_2063 : std_logic_vector(31 downto 0);
    signal call16_2066 : std_logic_vector(31 downto 0);
    signal call19_2069 : std_logic_vector(31 downto 0);
    signal call1_2051 : std_logic_vector(31 downto 0);
    signal call21_2072 : std_logic_vector(31 downto 0);
    signal call23_2075 : std_logic_vector(31 downto 0);
    signal call24_2078 : std_logic_vector(31 downto 0);
    signal call27_2081 : std_logic_vector(31 downto 0);
    signal call30_2084 : std_logic_vector(31 downto 0);
    signal call4_2054 : std_logic_vector(31 downto 0);
    signal call7_2057 : std_logic_vector(31 downto 0);
    signal call_2048 : std_logic_vector(31 downto 0);
    signal cmp112_2358 : std_logic_vector(0 downto 0);
    signal cmp128_2383 : std_logic_vector(0 downto 0);
    signal cmp_2328 : std_logic_vector(0 downto 0);
    signal conv100_2147 : std_logic_vector(31 downto 0);
    signal conv108_2353 : std_logic_vector(31 downto 0);
    signal conv111_2153 : std_logic_vector(31 downto 0);
    signal conv118_2378 : std_logic_vector(31 downto 0);
    signal conv121_2159 : std_logic_vector(31 downto 0);
    signal conv34_2091 : std_logic_vector(31 downto 0);
    signal conv35_2101 : std_logic_vector(15 downto 0);
    signal conv46_2215 : std_logic_vector(31 downto 0);
    signal conv48_2107 : std_logic_vector(31 downto 0);
    signal conv57_2229 : std_logic_vector(31 downto 0);
    signal conv71_2243 : std_logic_vector(31 downto 0);
    signal conv74_2135 : std_logic_vector(31 downto 0);
    signal conv76_2249 : std_logic_vector(31 downto 0);
    signal conv79_2141 : std_logic_vector(31 downto 0);
    signal conv81_2255 : std_logic_vector(31 downto 0);
    signal idxprom92_2306 : std_logic_vector(63 downto 0);
    signal idxprom_2285 : std_logic_vector(63 downto 0);
    signal inc116_2362 : std_logic_vector(15 downto 0);
    signal inc116x_xinput_dim0x_x2_2367 : std_logic_vector(15 downto 0);
    signal inc_2349 : std_logic_vector(15 downto 0);
    signal indvar_2173 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2416 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2404 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2194 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2398 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2187 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2374 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2391 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2180 : std_logic_vector(15 downto 0);
    signal mul60_2234 : std_logic_vector(31 downto 0);
    signal mul82_2260 : std_logic_vector(31 downto 0);
    signal mul84_2270 : std_logic_vector(31 downto 0);
    signal mul_2220 : std_logic_vector(31 downto 0);
    signal ptr_deref_2295_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2295_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2295_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2295_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2295_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2315_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2315_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2315_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2315_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2315_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2315_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr122143_2165 : std_logic_vector(31 downto 0);
    signal shr142_2097 : std_logic_vector(31 downto 0);
    signal shr87_2281 : std_logic_vector(31 downto 0);
    signal shr91_2302 : std_logic_vector(31 downto 0);
    signal sub54_2225 : std_logic_vector(31 downto 0);
    signal sub67_2129 : std_logic_vector(31 downto 0);
    signal sub68_2239 : std_logic_vector(31 downto 0);
    signal sub_2118 : std_logic_vector(31 downto 0);
    signal tmp1_2206 : std_logic_vector(31 downto 0);
    signal tmp89_2296 : std_logic_vector(63 downto 0);
    signal type_cast_2089_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2095_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2105_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2111_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2122_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2133_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2139_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2145_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2151_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2157_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2163_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2177_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2179_wire : std_logic_vector(31 downto 0);
    signal type_cast_2184_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2186_wire : std_logic_vector(15 downto 0);
    signal type_cast_2190_wire : std_logic_vector(15 downto 0);
    signal type_cast_2193_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2197_wire : std_logic_vector(15 downto 0);
    signal type_cast_2199_wire : std_logic_vector(15 downto 0);
    signal type_cast_2204_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2247_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2253_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2279_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2300_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2321_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2339_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2347_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2371_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2395_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2397_wire : std_logic_vector(15 downto 0);
    signal type_cast_2401_wire : std_logic_vector(15 downto 0);
    signal type_cast_2403_wire : std_logic_vector(15 downto 0);
    signal type_cast_2407_wire : std_logic_vector(15 downto 0);
    signal type_cast_2409_wire : std_logic_vector(15 downto 0);
    signal type_cast_2414_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2422_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_2290_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2290_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2290_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2290_resized_base_address <= "00000000000000";
    array_obj_ref_2311_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2311_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2311_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2311_resized_base_address <= "00000000000000";
    ptr_deref_2295_word_offset_0 <= "00000000000000";
    ptr_deref_2315_word_offset_0 <= "00000000000000";
    type_cast_2089_wire_constant <= "00000000000000000000000000000001";
    type_cast_2095_wire_constant <= "00000000000000000111111111111111";
    type_cast_2105_wire_constant <= "00000000000000001111111111111111";
    type_cast_2111_wire_constant <= "00000000000000001111111111111111";
    type_cast_2122_wire_constant <= "00000000000000001111111111111111";
    type_cast_2133_wire_constant <= "00000000000000001111111111111111";
    type_cast_2139_wire_constant <= "00000000000000001111111111111111";
    type_cast_2145_wire_constant <= "00000000000000001111111111111111";
    type_cast_2151_wire_constant <= "00000000000000001111111111111111";
    type_cast_2157_wire_constant <= "00000000000000000000000000000010";
    type_cast_2163_wire_constant <= "00000000000000000011111111111111";
    type_cast_2177_wire_constant <= "00000000000000000000000000000000";
    type_cast_2184_wire_constant <= "0000000000000000";
    type_cast_2193_wire_constant <= "0000000000000000";
    type_cast_2204_wire_constant <= "00000000000000000000000000000100";
    type_cast_2247_wire_constant <= "00000000000000001111111111111111";
    type_cast_2253_wire_constant <= "00000000000000001111111111111111";
    type_cast_2279_wire_constant <= "00000000000000000000000000000010";
    type_cast_2300_wire_constant <= "00000000000000000000000000000010";
    type_cast_2321_wire_constant <= "00000000000000000000000000000100";
    type_cast_2339_wire_constant <= "0000000000000100";
    type_cast_2347_wire_constant <= "0000000000000001";
    type_cast_2371_wire_constant <= "0000000000000000";
    type_cast_2395_wire_constant <= "0000000000000000";
    type_cast_2414_wire_constant <= "00000000000000000000000000000001";
    type_cast_2422_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_2173: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2177_wire_constant & type_cast_2179_wire;
      req <= phi_stmt_2173_req_0 & phi_stmt_2173_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2173",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2173_ack_0,
          idata => idata,
          odata => indvar_2173,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2173
    phi_stmt_2180: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2184_wire_constant & type_cast_2186_wire;
      req <= phi_stmt_2180_req_0 & phi_stmt_2180_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2180",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2180_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2180,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2180
    phi_stmt_2187: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2190_wire & type_cast_2193_wire_constant;
      req <= phi_stmt_2187_req_0 & phi_stmt_2187_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2187",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2187_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2187,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2187
    phi_stmt_2194: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2197_wire & type_cast_2199_wire;
      req <= phi_stmt_2194_req_0 & phi_stmt_2194_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2194",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2194_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2194,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2194
    phi_stmt_2391: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2395_wire_constant & type_cast_2397_wire;
      req <= phi_stmt_2391_req_0 & phi_stmt_2391_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2391",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2391_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2391,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2391
    phi_stmt_2398: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2401_wire & type_cast_2403_wire;
      req <= phi_stmt_2398_req_0 & phi_stmt_2398_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2398",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2398_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2398,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2398
    phi_stmt_2404: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2407_wire & type_cast_2409_wire;
      req <= phi_stmt_2404_req_0 & phi_stmt_2404_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2404",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2404_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2404,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2404
    -- flow-through select operator MUX_2373_inst
    input_dim1x_x2_2374 <= type_cast_2371_wire_constant when (cmp112_2358(0) /=  '0') else inc_2349;
    addr_of_2291_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2291_final_reg_req_0;
      addr_of_2291_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2291_final_reg_req_1;
      addr_of_2291_final_reg_ack_1<= rack(0);
      addr_of_2291_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2291_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2290_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx88_2292,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2312_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2312_final_reg_req_0;
      addr_of_2312_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2312_final_reg_req_1;
      addr_of_2312_final_reg_ack_1<= rack(0);
      addr_of_2312_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2312_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2311_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx93_2313,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2100_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2100_inst_req_0;
      type_cast_2100_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2100_inst_req_1;
      type_cast_2100_inst_ack_1<= rack(0);
      type_cast_2100_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2100_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr142_2097,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_2101,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2179_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2179_inst_req_0;
      type_cast_2179_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2179_inst_req_1;
      type_cast_2179_inst_ack_1<= rack(0);
      type_cast_2179_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2179_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2416,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2179_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2186_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2186_inst_req_0;
      type_cast_2186_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2186_inst_req_1;
      type_cast_2186_inst_ack_1<= rack(0);
      type_cast_2186_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2186_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2391,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2186_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2190_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2190_inst_req_0;
      type_cast_2190_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2190_inst_req_1;
      type_cast_2190_inst_ack_1<= rack(0);
      type_cast_2190_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2190_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2398,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2190_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2197_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2197_inst_req_0;
      type_cast_2197_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2197_inst_req_1;
      type_cast_2197_inst_ack_1<= rack(0);
      type_cast_2197_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2197_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv35_2101,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2197_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2199_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2199_inst_req_0;
      type_cast_2199_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2199_inst_req_1;
      type_cast_2199_inst_ack_1<= rack(0);
      type_cast_2199_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2199_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2404,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2199_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2214_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2214_inst_req_0;
      type_cast_2214_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2214_inst_req_1;
      type_cast_2214_inst_ack_1<= rack(0);
      type_cast_2214_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2214_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv46_2215,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2228_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2228_inst_req_0;
      type_cast_2228_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2228_inst_req_1;
      type_cast_2228_inst_ack_1<= rack(0);
      type_cast_2228_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2228_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2187,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv57_2229,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2242_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2242_inst_req_0;
      type_cast_2242_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2242_inst_req_1;
      type_cast_2242_inst_ack_1<= rack(0);
      type_cast_2242_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2242_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2180,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_2243,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2284_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2284_inst_req_0;
      type_cast_2284_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2284_inst_req_1;
      type_cast_2284_inst_ack_1<= rack(0);
      type_cast_2284_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2284_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr87_2281,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2285,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2305_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2305_inst_req_0;
      type_cast_2305_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2305_inst_req_1;
      type_cast_2305_inst_ack_1<= rack(0);
      type_cast_2305_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2305_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr91_2302,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom92_2306,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2352_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2352_inst_req_0;
      type_cast_2352_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2352_inst_req_1;
      type_cast_2352_inst_ack_1<= rack(0);
      type_cast_2352_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2352_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_2349,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv108_2353,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2361_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2361_inst_req_0;
      type_cast_2361_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2361_inst_req_1;
      type_cast_2361_inst_ack_1<= rack(0);
      type_cast_2361_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2361_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp112_2358,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc116_2362,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2377_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2377_inst_req_0;
      type_cast_2377_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2377_inst_req_1;
      type_cast_2377_inst_ack_1<= rack(0);
      type_cast_2377_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2377_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc116x_xinput_dim0x_x2_2367,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv118_2378,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2397_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2397_inst_req_0;
      type_cast_2397_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2397_inst_req_1;
      type_cast_2397_inst_ack_1<= rack(0);
      type_cast_2397_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2397_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add104_2341,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2397_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2401_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2401_inst_req_0;
      type_cast_2401_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2401_inst_req_1;
      type_cast_2401_inst_ack_1<= rack(0);
      type_cast_2401_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2401_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2374,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2401_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2403_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2403_inst_req_0;
      type_cast_2403_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2403_inst_req_1;
      type_cast_2403_inst_ack_1<= rack(0);
      type_cast_2403_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2403_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2187,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2403_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2407_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2407_inst_req_0;
      type_cast_2407_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2407_inst_req_1;
      type_cast_2407_inst_ack_1<= rack(0);
      type_cast_2407_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2407_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc116x_xinput_dim0x_x2_2367,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2407_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2409_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2409_inst_req_0;
      type_cast_2409_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2409_inst_req_1;
      type_cast_2409_inst_ack_1<= rack(0);
      type_cast_2409_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2409_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2409_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2290_index_1_rename
    process(R_idxprom_2289_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2289_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2289_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2290_index_1_resize
    process(idxprom_2285) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2285;
      ov := iv(13 downto 0);
      R_idxprom_2289_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2290_root_address_inst
    process(array_obj_ref_2290_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2290_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2290_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2311_index_1_rename
    process(R_idxprom92_2310_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom92_2310_resized;
      ov(13 downto 0) := iv;
      R_idxprom92_2310_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2311_index_1_resize
    process(idxprom92_2306) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom92_2306;
      ov := iv(13 downto 0);
      R_idxprom92_2310_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2311_root_address_inst
    process(array_obj_ref_2311_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2311_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2311_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2295_addr_0
    process(ptr_deref_2295_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2295_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2295_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2295_base_resize
    process(arrayidx88_2292) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx88_2292;
      ov := iv(13 downto 0);
      ptr_deref_2295_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2295_gather_scatter
    process(ptr_deref_2295_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2295_data_0;
      ov(63 downto 0) := iv;
      tmp89_2296 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2295_root_address_inst
    process(ptr_deref_2295_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2295_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2295_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2315_addr_0
    process(ptr_deref_2315_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2315_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2315_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2315_base_resize
    process(arrayidx93_2313) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx93_2313;
      ov := iv(13 downto 0);
      ptr_deref_2315_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2315_gather_scatter
    process(tmp89_2296) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp89_2296;
      ov(63 downto 0) := iv;
      ptr_deref_2315_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2315_root_address_inst
    process(ptr_deref_2315_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2315_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2315_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2329_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2328;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2329_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2329_branch_req_0,
          ack0 => if_stmt_2329_branch_ack_0,
          ack1 => if_stmt_2329_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2384_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp128_2383;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2384_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2384_branch_req_0,
          ack0 => if_stmt_2384_branch_ack_0,
          ack1 => if_stmt_2384_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2340_inst
    process(input_dim2x_x1_2180) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2180, type_cast_2339_wire_constant, tmp_var);
      add104_2341 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2348_inst
    process(input_dim1x_x1_2187) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2187, type_cast_2347_wire_constant, tmp_var);
      inc_2349 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2366_inst
    process(inc116_2362, input_dim0x_x2_2194) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc116_2362, input_dim0x_x2_2194, tmp_var);
      inc116x_xinput_dim0x_x2_2367 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2112_inst
    process(call10_2060) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call10_2060, type_cast_2111_wire_constant, tmp_var);
      add_2113 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2123_inst
    process(call13_2063) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call13_2063, type_cast_2122_wire_constant, tmp_var);
      add64_2124 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2169_inst
    process(shr122143_2165, shr142_2097) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr122143_2165, shr142_2097, tmp_var);
      add127_2170 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2210_inst
    process(call23_2075, tmp1_2206) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call23_2075, tmp1_2206, tmp_var);
      add_src_0x_x0_2211 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2224_inst
    process(sub_2118, mul_2220) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2118, mul_2220, tmp_var);
      sub54_2225 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2238_inst
    process(sub67_2129, mul60_2234) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub67_2129, mul60_2234, tmp_var);
      sub68_2239 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2264_inst
    process(mul82_2260, conv76_2249) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul82_2260, conv76_2249, tmp_var);
      add83_2265 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2274_inst
    process(mul84_2270, conv71_2243) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul84_2270, conv71_2243, tmp_var);
      add85_2275 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2322_inst
    process(conv71_2243) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv71_2243, type_cast_2321_wire_constant, tmp_var);
      add97_2323 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2415_inst
    process(indvar_2173) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2173, type_cast_2414_wire_constant, tmp_var);
      indvarx_xnext_2416 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2096_inst
    process(conv34_2091) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv34_2091, type_cast_2095_wire_constant, tmp_var);
      shr142_2097 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2106_inst
    process(call19_2069) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call19_2069, type_cast_2105_wire_constant, tmp_var);
      conv48_2107 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2134_inst
    process(call30_2084) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call30_2084, type_cast_2133_wire_constant, tmp_var);
      conv74_2135 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2140_inst
    process(call27_2081) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call27_2081, type_cast_2139_wire_constant, tmp_var);
      conv79_2141 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2146_inst
    process(call4_2054) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call4_2054, type_cast_2145_wire_constant, tmp_var);
      conv100_2147 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2152_inst
    process(call1_2051) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call1_2051, type_cast_2151_wire_constant, tmp_var);
      conv111_2153 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2164_inst
    process(conv121_2159) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv121_2159, type_cast_2163_wire_constant, tmp_var);
      shr122143_2165 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2248_inst
    process(sub68_2239) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(sub68_2239, type_cast_2247_wire_constant, tmp_var);
      conv76_2249 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2254_inst
    process(sub54_2225) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(sub54_2225, type_cast_2253_wire_constant, tmp_var);
      conv81_2255 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2357_inst
    process(conv108_2353, conv111_2153) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv108_2353, conv111_2153, tmp_var);
      cmp112_2358 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2382_inst
    process(conv118_2378, add127_2170) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv118_2378, add127_2170, tmp_var);
      cmp128_2383 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2090_inst
    process(call_2048) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2048, type_cast_2089_wire_constant, tmp_var);
      conv34_2091 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2158_inst
    process(call_2048) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2048, type_cast_2157_wire_constant, tmp_var);
      conv121_2159 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2280_inst
    process(add_src_0x_x0_2211) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2211, type_cast_2279_wire_constant, tmp_var);
      shr87_2281 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2301_inst
    process(add85_2275) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add85_2275, type_cast_2300_wire_constant, tmp_var);
      shr91_2302 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2205_inst
    process(indvar_2173) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2173, type_cast_2204_wire_constant, tmp_var);
      tmp1_2206 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2219_inst
    process(conv46_2215, conv48_2107) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv46_2215, conv48_2107, tmp_var);
      mul_2220 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2233_inst
    process(conv57_2229, conv48_2107) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv57_2229, conv48_2107, tmp_var);
      mul60_2234 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2259_inst
    process(conv81_2255, conv79_2141) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv81_2255, conv79_2141, tmp_var);
      mul82_2260 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2269_inst
    process(add83_2265, conv74_2135) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add83_2265, conv74_2135, tmp_var);
      mul84_2270 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2117_inst
    process(add_2113, call21_2072) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add_2113, call21_2072, tmp_var);
      sub_2118 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2128_inst
    process(add64_2124, call21_2072) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add64_2124, call21_2072, tmp_var);
      sub67_2129 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2327_inst
    process(add97_2323, conv100_2147) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add97_2323, conv100_2147, tmp_var);
      cmp_2328 <= tmp_var; --
    end process;
    -- shared split operator group (36) : array_obj_ref_2290_index_offset 
    ApIntAdd_group_36: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2289_scaled;
      array_obj_ref_2290_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2290_index_offset_req_0;
      array_obj_ref_2290_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2290_index_offset_req_1;
      array_obj_ref_2290_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_36_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : array_obj_ref_2311_index_offset 
    ApIntAdd_group_37: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom92_2310_scaled;
      array_obj_ref_2311_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2311_index_offset_req_0;
      array_obj_ref_2311_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2311_index_offset_req_1;
      array_obj_ref_2311_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_37_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_37_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_37",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared load operator group (0) : ptr_deref_2295_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2295_load_0_req_0;
      ptr_deref_2295_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2295_load_0_req_1;
      ptr_deref_2295_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2295_word_address_0;
      ptr_deref_2295_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2315_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2315_store_0_req_0;
      ptr_deref_2315_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2315_store_0_req_1;
      ptr_deref_2315_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2315_word_address_0;
      data_in <= ptr_deref_2315_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2047_inst RPIPE_Block2_start_2050_inst RPIPE_Block2_start_2053_inst RPIPE_Block2_start_2056_inst RPIPE_Block2_start_2059_inst RPIPE_Block2_start_2062_inst RPIPE_Block2_start_2065_inst RPIPE_Block2_start_2068_inst RPIPE_Block2_start_2071_inst RPIPE_Block2_start_2074_inst RPIPE_Block2_start_2077_inst RPIPE_Block2_start_2080_inst RPIPE_Block2_start_2083_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(415 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 12 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 12 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 12 downto 0);
      signal guard_vector : std_logic_vector( 12 downto 0);
      constant outBUFs : IntegerArray(12 downto 0) := (12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(12 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false);
      constant guardBuffering: IntegerArray(12 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2);
      -- 
    begin -- 
      reqL_unguarded(12) <= RPIPE_Block2_start_2047_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block2_start_2050_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block2_start_2053_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block2_start_2056_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block2_start_2059_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block2_start_2062_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block2_start_2065_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block2_start_2068_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block2_start_2071_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block2_start_2074_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block2_start_2077_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block2_start_2080_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block2_start_2083_inst_req_0;
      RPIPE_Block2_start_2047_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block2_start_2050_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block2_start_2053_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block2_start_2056_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block2_start_2059_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block2_start_2062_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block2_start_2065_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block2_start_2068_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block2_start_2071_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block2_start_2074_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block2_start_2077_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block2_start_2080_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block2_start_2083_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(12) <= RPIPE_Block2_start_2047_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block2_start_2050_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block2_start_2053_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block2_start_2056_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block2_start_2059_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block2_start_2062_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block2_start_2065_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block2_start_2068_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block2_start_2071_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block2_start_2074_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block2_start_2077_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block2_start_2080_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block2_start_2083_inst_req_1;
      RPIPE_Block2_start_2047_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block2_start_2050_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block2_start_2053_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block2_start_2056_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block2_start_2059_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block2_start_2062_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block2_start_2065_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block2_start_2068_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block2_start_2071_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block2_start_2074_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block2_start_2077_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block2_start_2080_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block2_start_2083_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      call_2048 <= data_out(415 downto 384);
      call1_2051 <= data_out(383 downto 352);
      call4_2054 <= data_out(351 downto 320);
      call7_2057 <= data_out(319 downto 288);
      call10_2060 <= data_out(287 downto 256);
      call13_2063 <= data_out(255 downto 224);
      call16_2066 <= data_out(223 downto 192);
      call19_2069 <= data_out(191 downto 160);
      call21_2072 <= data_out(159 downto 128);
      call23_2075 <= data_out(127 downto 96);
      call24_2078 <= data_out(95 downto 64);
      call27_2081 <= data_out(63 downto 32);
      call30_2084 <= data_out(31 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 13, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 32,  num_reqs => 13,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2420_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2420_inst_req_0;
      WPIPE_Block2_done_2420_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2420_inst_req_1;
      WPIPE_Block2_done_2420_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2422_wire_constant;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(31 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_6059_start: Boolean;
  signal convTransposeD_CP_6059_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal addr_of_2702_final_reg_req_1 : boolean;
  signal type_cast_2767_inst_ack_1 : boolean;
  signal ptr_deref_2705_store_0_ack_1 : boolean;
  signal type_cast_2742_inst_ack_1 : boolean;
  signal ptr_deref_2705_store_0_req_0 : boolean;
  signal ptr_deref_2705_store_0_req_1 : boolean;
  signal type_cast_2751_inst_req_1 : boolean;
  signal addr_of_2702_final_reg_ack_0 : boolean;
  signal addr_of_2702_final_reg_req_0 : boolean;
  signal type_cast_2751_inst_ack_1 : boolean;
  signal type_cast_2767_inst_req_0 : boolean;
  signal if_stmt_2719_branch_ack_0 : boolean;
  signal ptr_deref_2705_store_0_ack_0 : boolean;
  signal addr_of_2702_final_reg_ack_1 : boolean;
  signal type_cast_2767_inst_req_1 : boolean;
  signal WPIPE_Block3_done_2810_inst_req_1 : boolean;
  signal phi_stmt_2570_req_1 : boolean;
  signal WPIPE_Block3_done_2810_inst_ack_1 : boolean;
  signal type_cast_2767_inst_ack_0 : boolean;
  signal if_stmt_2719_branch_req_0 : boolean;
  signal type_cast_2587_inst_req_1 : boolean;
  signal type_cast_2587_inst_ack_1 : boolean;
  signal phi_stmt_2563_req_1 : boolean;
  signal type_cast_2751_inst_req_0 : boolean;
  signal type_cast_2751_inst_ack_0 : boolean;
  signal if_stmt_2719_branch_ack_1 : boolean;
  signal phi_stmt_2577_req_1 : boolean;
  signal type_cast_2587_inst_req_0 : boolean;
  signal phi_stmt_2584_req_0 : boolean;
  signal type_cast_2587_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2431_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2431_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2431_inst_req_1 : boolean;
  signal type_cast_2742_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2431_inst_ack_1 : boolean;
  signal WPIPE_Block3_done_2810_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_2810_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2434_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2434_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2434_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2434_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2437_inst_req_0 : boolean;
  signal type_cast_2742_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2437_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2437_inst_req_1 : boolean;
  signal type_cast_2742_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2437_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2440_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2440_inst_ack_0 : boolean;
  signal array_obj_ref_2701_index_offset_ack_1 : boolean;
  signal RPIPE_Block3_start_2440_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2440_inst_ack_1 : boolean;
  signal array_obj_ref_2701_index_offset_req_1 : boolean;
  signal if_stmt_2774_branch_ack_0 : boolean;
  signal if_stmt_2774_branch_ack_1 : boolean;
  signal RPIPE_Block3_start_2443_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2443_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2443_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2443_inst_ack_1 : boolean;
  signal if_stmt_2774_branch_req_0 : boolean;
  signal RPIPE_Block3_start_2446_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2446_inst_ack_0 : boolean;
  signal array_obj_ref_2701_index_offset_ack_0 : boolean;
  signal RPIPE_Block3_start_2446_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2446_inst_ack_1 : boolean;
  signal array_obj_ref_2701_index_offset_req_0 : boolean;
  signal RPIPE_Block3_start_2449_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2449_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2449_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2449_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2452_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2452_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2452_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2452_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2455_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2455_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2455_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2455_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2458_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2458_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2458_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2458_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2461_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2461_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2461_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2461_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2464_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2464_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2464_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2464_inst_ack_1 : boolean;
  signal RPIPE_Block3_start_2467_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2467_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2467_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2467_inst_ack_1 : boolean;
  signal type_cast_2501_inst_req_0 : boolean;
  signal type_cast_2501_inst_ack_0 : boolean;
  signal type_cast_2501_inst_req_1 : boolean;
  signal type_cast_2501_inst_ack_1 : boolean;
  signal type_cast_2604_inst_req_0 : boolean;
  signal type_cast_2604_inst_ack_0 : boolean;
  signal type_cast_2604_inst_req_1 : boolean;
  signal type_cast_2604_inst_ack_1 : boolean;
  signal type_cast_2618_inst_req_0 : boolean;
  signal type_cast_2618_inst_ack_0 : boolean;
  signal type_cast_2618_inst_req_1 : boolean;
  signal type_cast_2618_inst_ack_1 : boolean;
  signal type_cast_2632_inst_req_0 : boolean;
  signal type_cast_2632_inst_ack_0 : boolean;
  signal type_cast_2632_inst_req_1 : boolean;
  signal type_cast_2632_inst_ack_1 : boolean;
  signal type_cast_2674_inst_req_0 : boolean;
  signal type_cast_2674_inst_ack_0 : boolean;
  signal type_cast_2674_inst_req_1 : boolean;
  signal type_cast_2674_inst_ack_1 : boolean;
  signal array_obj_ref_2680_index_offset_req_0 : boolean;
  signal array_obj_ref_2680_index_offset_ack_0 : boolean;
  signal array_obj_ref_2680_index_offset_req_1 : boolean;
  signal array_obj_ref_2680_index_offset_ack_1 : boolean;
  signal addr_of_2681_final_reg_req_0 : boolean;
  signal addr_of_2681_final_reg_ack_0 : boolean;
  signal addr_of_2681_final_reg_req_1 : boolean;
  signal addr_of_2681_final_reg_ack_1 : boolean;
  signal ptr_deref_2685_load_0_req_0 : boolean;
  signal ptr_deref_2685_load_0_ack_0 : boolean;
  signal ptr_deref_2685_load_0_req_1 : boolean;
  signal ptr_deref_2685_load_0_ack_1 : boolean;
  signal type_cast_2695_inst_req_0 : boolean;
  signal type_cast_2695_inst_ack_0 : boolean;
  signal type_cast_2695_inst_req_1 : boolean;
  signal type_cast_2695_inst_ack_1 : boolean;
  signal type_cast_2566_inst_req_0 : boolean;
  signal type_cast_2566_inst_ack_0 : boolean;
  signal type_cast_2566_inst_req_1 : boolean;
  signal type_cast_2566_inst_ack_1 : boolean;
  signal phi_stmt_2563_req_0 : boolean;
  signal type_cast_2573_inst_req_0 : boolean;
  signal type_cast_2573_inst_ack_0 : boolean;
  signal type_cast_2573_inst_req_1 : boolean;
  signal type_cast_2573_inst_ack_1 : boolean;
  signal phi_stmt_2570_req_0 : boolean;
  signal type_cast_2580_inst_req_0 : boolean;
  signal type_cast_2580_inst_ack_0 : boolean;
  signal type_cast_2580_inst_req_1 : boolean;
  signal type_cast_2580_inst_ack_1 : boolean;
  signal phi_stmt_2577_req_0 : boolean;
  signal type_cast_2589_inst_req_0 : boolean;
  signal type_cast_2589_inst_ack_0 : boolean;
  signal type_cast_2589_inst_req_1 : boolean;
  signal type_cast_2589_inst_ack_1 : boolean;
  signal phi_stmt_2584_req_1 : boolean;
  signal phi_stmt_2563_ack_0 : boolean;
  signal phi_stmt_2570_ack_0 : boolean;
  signal phi_stmt_2577_ack_0 : boolean;
  signal phi_stmt_2584_ack_0 : boolean;
  signal phi_stmt_2781_req_1 : boolean;
  signal type_cast_2793_inst_req_0 : boolean;
  signal type_cast_2793_inst_ack_0 : boolean;
  signal type_cast_2793_inst_req_1 : boolean;
  signal type_cast_2793_inst_ack_1 : boolean;
  signal phi_stmt_2788_req_1 : boolean;
  signal type_cast_2799_inst_req_0 : boolean;
  signal type_cast_2799_inst_ack_0 : boolean;
  signal type_cast_2799_inst_req_1 : boolean;
  signal type_cast_2799_inst_ack_1 : boolean;
  signal phi_stmt_2794_req_1 : boolean;
  signal type_cast_2784_inst_req_0 : boolean;
  signal type_cast_2784_inst_ack_0 : boolean;
  signal type_cast_2784_inst_req_1 : boolean;
  signal type_cast_2784_inst_ack_1 : boolean;
  signal phi_stmt_2781_req_0 : boolean;
  signal type_cast_2791_inst_req_0 : boolean;
  signal type_cast_2791_inst_ack_0 : boolean;
  signal type_cast_2791_inst_req_1 : boolean;
  signal type_cast_2791_inst_ack_1 : boolean;
  signal phi_stmt_2788_req_0 : boolean;
  signal type_cast_2797_inst_req_0 : boolean;
  signal type_cast_2797_inst_ack_0 : boolean;
  signal type_cast_2797_inst_req_1 : boolean;
  signal type_cast_2797_inst_ack_1 : boolean;
  signal phi_stmt_2794_req_0 : boolean;
  signal phi_stmt_2781_ack_0 : boolean;
  signal phi_stmt_2788_ack_0 : boolean;
  signal phi_stmt_2794_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_6059_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6059_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_6059_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_6059_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_6059: Block -- control-path 
    signal convTransposeD_CP_6059_elements: BooleanArray(115 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_6059_elements(0) <= convTransposeD_CP_6059_start;
    convTransposeD_CP_6059_symbol <= convTransposeD_CP_6059_elements(66);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2429/branch_block_stmt_2429__entry__
      -- CP-element group 0: 	 branch_block_stmt_2429/$entry
      -- CP-element group 0: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/$entry
      -- CP-element group 0: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2431_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2431_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2431_Sample/rr
      -- 
    rr_6107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(0), ack => RPIPE_Block3_start_2431_inst_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	115 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	74 
    -- CP-element group 1: 	75 
    -- CP-element group 1: 	77 
    -- CP-element group 1: 	78 
    -- CP-element group 1: 	80 
    -- CP-element group 1: 	81 
    -- CP-element group 1: 	83 
    -- CP-element group 1: 	84 
    -- CP-element group 1:  members (39) 
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody
      -- CP-element group 1: 	 branch_block_stmt_2429/assign_stmt_2806__exit__
      -- CP-element group 1: 	 branch_block_stmt_2429/assign_stmt_2806__entry__
      -- CP-element group 1: 	 branch_block_stmt_2429/merge_stmt_2780__exit__
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2563/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/assign_stmt_2806/$exit
      -- CP-element group 1: 	 branch_block_stmt_2429/assign_stmt_2806/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2570/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_sources/type_cast_2573/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_sources/type_cast_2573/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_sources/type_cast_2573/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_sources/type_cast_2573/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_sources/type_cast_2573/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_sources/type_cast_2573/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2577/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_sources/type_cast_2580/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_sources/type_cast_2580/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_sources/type_cast_2580/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_sources/type_cast_2580/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_sources/type_cast_2580/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_sources/type_cast_2580/SplitProtocol/Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2584/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2589/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2589/SplitProtocol/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2589/SplitProtocol/Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2589/SplitProtocol/Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2589/SplitProtocol/Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2589/SplitProtocol/Update/cr
      -- 
    rr_6738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(1), ack => type_cast_2566_inst_req_0); -- 
    cr_6743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(1), ack => type_cast_2566_inst_req_1); -- 
    rr_6761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(1), ack => type_cast_2573_inst_req_0); -- 
    cr_6766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(1), ack => type_cast_2573_inst_req_1); -- 
    rr_6784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(1), ack => type_cast_2580_inst_req_0); -- 
    cr_6789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(1), ack => type_cast_2580_inst_req_1); -- 
    rr_6807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(1), ack => type_cast_2589_inst_req_0); -- 
    cr_6812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(1), ack => type_cast_2589_inst_req_1); -- 
    convTransposeD_CP_6059_elements(1) <= convTransposeD_CP_6059_elements(115);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2431_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2431_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2431_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2431_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2431_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2431_Update/cr
      -- 
    ra_6108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2431_inst_ack_0, ack => convTransposeD_CP_6059_elements(2)); -- 
    cr_6112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(2), ack => RPIPE_Block3_start_2431_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2431_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2431_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2431_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2434_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2434_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2434_Sample/rr
      -- 
    ca_6113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2431_inst_ack_1, ack => convTransposeD_CP_6059_elements(3)); -- 
    rr_6121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(3), ack => RPIPE_Block3_start_2434_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2434_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2434_update_start_
      -- CP-element group 4: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2434_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2434_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2434_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2434_Update/cr
      -- 
    ra_6122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2434_inst_ack_0, ack => convTransposeD_CP_6059_elements(4)); -- 
    cr_6126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(4), ack => RPIPE_Block3_start_2434_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2434_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2434_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2434_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2437_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2437_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2437_Sample/rr
      -- 
    ca_6127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2434_inst_ack_1, ack => convTransposeD_CP_6059_elements(5)); -- 
    rr_6135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(5), ack => RPIPE_Block3_start_2437_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2437_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2437_update_start_
      -- CP-element group 6: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2437_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2437_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2437_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2437_Update/cr
      -- 
    ra_6136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2437_inst_ack_0, ack => convTransposeD_CP_6059_elements(6)); -- 
    cr_6140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(6), ack => RPIPE_Block3_start_2437_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2437_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2437_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2437_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2440_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2440_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2440_Sample/rr
      -- 
    ca_6141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2437_inst_ack_1, ack => convTransposeD_CP_6059_elements(7)); -- 
    rr_6149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(7), ack => RPIPE_Block3_start_2440_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2440_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2440_update_start_
      -- CP-element group 8: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2440_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2440_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2440_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2440_Update/cr
      -- 
    ra_6150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2440_inst_ack_0, ack => convTransposeD_CP_6059_elements(8)); -- 
    cr_6154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(8), ack => RPIPE_Block3_start_2440_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2440_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2440_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2440_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2443_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2443_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2443_Sample/rr
      -- 
    ca_6155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2440_inst_ack_1, ack => convTransposeD_CP_6059_elements(9)); -- 
    rr_6163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(9), ack => RPIPE_Block3_start_2443_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2443_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2443_update_start_
      -- CP-element group 10: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2443_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2443_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2443_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2443_Update/cr
      -- 
    ra_6164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2443_inst_ack_0, ack => convTransposeD_CP_6059_elements(10)); -- 
    cr_6168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(10), ack => RPIPE_Block3_start_2443_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2443_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2443_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2443_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2446_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2446_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2446_Sample/rr
      -- 
    ca_6169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2443_inst_ack_1, ack => convTransposeD_CP_6059_elements(11)); -- 
    rr_6177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(11), ack => RPIPE_Block3_start_2446_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2446_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2446_update_start_
      -- CP-element group 12: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2446_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2446_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2446_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2446_Update/cr
      -- 
    ra_6178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2446_inst_ack_0, ack => convTransposeD_CP_6059_elements(12)); -- 
    cr_6182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(12), ack => RPIPE_Block3_start_2446_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2446_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2446_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2446_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2449_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2449_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2449_Sample/rr
      -- 
    ca_6183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2446_inst_ack_1, ack => convTransposeD_CP_6059_elements(13)); -- 
    rr_6191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(13), ack => RPIPE_Block3_start_2449_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2449_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2449_update_start_
      -- CP-element group 14: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2449_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2449_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2449_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2449_Update/cr
      -- 
    ra_6192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2449_inst_ack_0, ack => convTransposeD_CP_6059_elements(14)); -- 
    cr_6196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(14), ack => RPIPE_Block3_start_2449_inst_req_1); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2449_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2449_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2449_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2452_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2452_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2452_Sample/rr
      -- 
    ca_6197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2449_inst_ack_1, ack => convTransposeD_CP_6059_elements(15)); -- 
    rr_6205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(15), ack => RPIPE_Block3_start_2452_inst_req_0); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (6) 
      -- CP-element group 16: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2452_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2452_update_start_
      -- CP-element group 16: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2452_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2452_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2452_Update/$entry
      -- CP-element group 16: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2452_Update/cr
      -- 
    ra_6206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2452_inst_ack_0, ack => convTransposeD_CP_6059_elements(16)); -- 
    cr_6210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(16), ack => RPIPE_Block3_start_2452_inst_req_1); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2452_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2452_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2452_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2455_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2455_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2455_Sample/rr
      -- 
    ca_6211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2452_inst_ack_1, ack => convTransposeD_CP_6059_elements(17)); -- 
    rr_6219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(17), ack => RPIPE_Block3_start_2455_inst_req_0); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2455_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2455_update_start_
      -- CP-element group 18: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2455_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2455_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2455_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2455_Update/cr
      -- 
    ra_6220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2455_inst_ack_0, ack => convTransposeD_CP_6059_elements(18)); -- 
    cr_6224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(18), ack => RPIPE_Block3_start_2455_inst_req_1); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2455_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2455_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2455_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2458_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2458_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2458_Sample/rr
      -- 
    ca_6225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2455_inst_ack_1, ack => convTransposeD_CP_6059_elements(19)); -- 
    rr_6233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(19), ack => RPIPE_Block3_start_2458_inst_req_0); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (6) 
      -- CP-element group 20: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2458_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2458_update_start_
      -- CP-element group 20: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2458_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2458_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2458_Update/$entry
      -- CP-element group 20: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2458_Update/cr
      -- 
    ra_6234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2458_inst_ack_0, ack => convTransposeD_CP_6059_elements(20)); -- 
    cr_6238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(20), ack => RPIPE_Block3_start_2458_inst_req_1); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2458_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2458_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2458_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2461_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2461_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2461_Sample/rr
      -- 
    ca_6239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2458_inst_ack_1, ack => convTransposeD_CP_6059_elements(21)); -- 
    rr_6247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(21), ack => RPIPE_Block3_start_2461_inst_req_0); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2461_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2461_update_start_
      -- CP-element group 22: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2461_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2461_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2461_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2461_Update/cr
      -- 
    ra_6248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2461_inst_ack_0, ack => convTransposeD_CP_6059_elements(22)); -- 
    cr_6252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(22), ack => RPIPE_Block3_start_2461_inst_req_1); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2461_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2461_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2461_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2464_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2464_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2464_Sample/rr
      -- 
    ca_6253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2461_inst_ack_1, ack => convTransposeD_CP_6059_elements(23)); -- 
    rr_6261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(23), ack => RPIPE_Block3_start_2464_inst_req_0); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2464_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2464_update_start_
      -- CP-element group 24: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2464_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2464_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2464_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2464_Update/cr
      -- 
    ra_6262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2464_inst_ack_0, ack => convTransposeD_CP_6059_elements(24)); -- 
    cr_6266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(24), ack => RPIPE_Block3_start_2464_inst_req_1); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2464_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2464_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2464_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2467_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2467_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2467_Sample/rr
      -- 
    ca_6267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2464_inst_ack_1, ack => convTransposeD_CP_6059_elements(25)); -- 
    rr_6275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(25), ack => RPIPE_Block3_start_2467_inst_req_0); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2467_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2467_update_start_
      -- CP-element group 26: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2467_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2467_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2467_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2467_Update/cr
      -- 
    ra_6276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2467_inst_ack_0, ack => convTransposeD_CP_6059_elements(26)); -- 
    cr_6280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(26), ack => RPIPE_Block3_start_2467_inst_req_1); -- 
    -- CP-element group 27:  fork  transition  place  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (13) 
      -- CP-element group 27: 	 branch_block_stmt_2429/assign_stmt_2475_to_assign_stmt_2560__entry__
      -- CP-element group 27: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468__exit__
      -- CP-element group 27: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/$exit
      -- CP-element group 27: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2467_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2467_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_2429/assign_stmt_2432_to_assign_stmt_2468/RPIPE_Block3_start_2467_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_2429/assign_stmt_2475_to_assign_stmt_2560/$entry
      -- CP-element group 27: 	 branch_block_stmt_2429/assign_stmt_2475_to_assign_stmt_2560/type_cast_2501_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_2429/assign_stmt_2475_to_assign_stmt_2560/type_cast_2501_update_start_
      -- CP-element group 27: 	 branch_block_stmt_2429/assign_stmt_2475_to_assign_stmt_2560/type_cast_2501_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_2429/assign_stmt_2475_to_assign_stmt_2560/type_cast_2501_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_2429/assign_stmt_2475_to_assign_stmt_2560/type_cast_2501_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_2429/assign_stmt_2475_to_assign_stmt_2560/type_cast_2501_Update/cr
      -- 
    ca_6281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2467_inst_ack_1, ack => convTransposeD_CP_6059_elements(27)); -- 
    rr_6292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(27), ack => type_cast_2501_inst_req_0); -- 
    cr_6297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(27), ack => type_cast_2501_inst_req_1); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2429/assign_stmt_2475_to_assign_stmt_2560/type_cast_2501_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_2429/assign_stmt_2475_to_assign_stmt_2560/type_cast_2501_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_2429/assign_stmt_2475_to_assign_stmt_2560/type_cast_2501_Sample/ra
      -- 
    ra_6293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2501_inst_ack_0, ack => convTransposeD_CP_6059_elements(28)); -- 
    -- CP-element group 29:  fork  transition  place  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	67 
    -- CP-element group 29: 	68 
    -- CP-element group 29: 	69 
    -- CP-element group 29: 	70 
    -- CP-element group 29: 	71 
    -- CP-element group 29:  members (21) 
      -- CP-element group 29: 	 branch_block_stmt_2429/entry_whilex_xbody
      -- CP-element group 29: 	 branch_block_stmt_2429/assign_stmt_2475_to_assign_stmt_2560__exit__
      -- CP-element group 29: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2587/SplitProtocol/Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2587/SplitProtocol/Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2584/$entry
      -- CP-element group 29: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2570/$entry
      -- CP-element group 29: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2587/SplitProtocol/Update/cr
      -- CP-element group 29: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2587/$entry
      -- CP-element group 29: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/$entry
      -- CP-element group 29: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2563/$entry
      -- CP-element group 29: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2577/$entry
      -- CP-element group 29: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2587/SplitProtocol/$entry
      -- CP-element group 29: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2587/SplitProtocol/Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_2429/assign_stmt_2475_to_assign_stmt_2560/$exit
      -- CP-element group 29: 	 branch_block_stmt_2429/assign_stmt_2475_to_assign_stmt_2560/type_cast_2501_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_2429/assign_stmt_2475_to_assign_stmt_2560/type_cast_2501_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_2429/assign_stmt_2475_to_assign_stmt_2560/type_cast_2501_Update/ca
      -- 
    ca_6298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2501_inst_ack_1, ack => convTransposeD_CP_6059_elements(29)); -- 
    cr_6717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(29), ack => type_cast_2587_inst_req_1); -- 
    rr_6712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(29), ack => type_cast_2587_inst_req_0); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	92 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2604_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2604_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2604_Sample/ra
      -- 
    ra_6310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2604_inst_ack_0, ack => convTransposeD_CP_6059_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	92 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	44 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2604_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2604_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2604_Update/ca
      -- 
    ca_6315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2604_inst_ack_1, ack => convTransposeD_CP_6059_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	92 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2618_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2618_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2618_Sample/ra
      -- 
    ra_6324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2618_inst_ack_0, ack => convTransposeD_CP_6059_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	92 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	44 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2618_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2618_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2618_Update/ca
      -- 
    ca_6329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2618_inst_ack_1, ack => convTransposeD_CP_6059_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	92 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2632_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2632_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2632_Sample/ra
      -- 
    ra_6338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2632_inst_ack_0, ack => convTransposeD_CP_6059_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	92 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	44 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2632_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2632_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2632_Update/ca
      -- 
    ca_6343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2632_inst_ack_1, ack => convTransposeD_CP_6059_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	92 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2674_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2674_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2674_Sample/ra
      -- 
    ra_6352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2674_inst_ack_0, ack => convTransposeD_CP_6059_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	92 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (16) 
      -- CP-element group 37: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2674_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2674_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2674_Update/ca
      -- CP-element group 37: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_index_resized_1
      -- CP-element group 37: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_index_scaled_1
      -- CP-element group 37: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_index_computed_1
      -- CP-element group 37: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_index_resize_1/$entry
      -- CP-element group 37: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_index_resize_1/$exit
      -- CP-element group 37: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_index_resize_1/index_resize_req
      -- CP-element group 37: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_index_resize_1/index_resize_ack
      -- CP-element group 37: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_index_scale_1/$entry
      -- CP-element group 37: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_index_scale_1/$exit
      -- CP-element group 37: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_index_scale_1/scale_rename_req
      -- CP-element group 37: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_index_scale_1/scale_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_final_index_sum_regn_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_final_index_sum_regn_Sample/req
      -- 
    ca_6357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2674_inst_ack_1, ack => convTransposeD_CP_6059_elements(37)); -- 
    req_6382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(37), ack => array_obj_ref_2680_index_offset_req_0); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	54 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_final_index_sum_regn_sample_complete
      -- CP-element group 38: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_final_index_sum_regn_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_final_index_sum_regn_Sample/ack
      -- 
    ack_6383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2680_index_offset_ack_0, ack => convTransposeD_CP_6059_elements(38)); -- 
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	92 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (11) 
      -- CP-element group 39: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2681_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_root_address_calculated
      -- CP-element group 39: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_offset_calculated
      -- CP-element group 39: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_final_index_sum_regn_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_final_index_sum_regn_Update/ack
      -- CP-element group 39: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_base_plus_offset/$entry
      -- CP-element group 39: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_base_plus_offset/$exit
      -- CP-element group 39: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_base_plus_offset/sum_rename_req
      -- CP-element group 39: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_base_plus_offset/sum_rename_ack
      -- CP-element group 39: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2681_request/$entry
      -- CP-element group 39: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2681_request/req
      -- 
    ack_6388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2680_index_offset_ack_1, ack => convTransposeD_CP_6059_elements(39)); -- 
    req_6397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(39), ack => addr_of_2681_final_reg_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2681_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2681_request/$exit
      -- CP-element group 40: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2681_request/ack
      -- 
    ack_6398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2681_final_reg_ack_0, ack => convTransposeD_CP_6059_elements(40)); -- 
    -- CP-element group 41:  join  fork  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	92 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (24) 
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2681_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2681_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2681_complete/ack
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_base_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_word_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_base_address_resized
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_base_addr_resize/$entry
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_base_addr_resize/$exit
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_base_addr_resize/base_resize_req
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_base_addr_resize/base_resize_ack
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_base_plus_offset/$entry
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_base_plus_offset/$exit
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_word_addrgen/$entry
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_word_addrgen/$exit
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_word_addrgen/root_register_req
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_word_addrgen/root_register_ack
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Sample/word_access_start/$entry
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Sample/word_access_start/word_0/$entry
      -- CP-element group 41: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Sample/word_access_start/word_0/rr
      -- 
    ack_6403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2681_final_reg_ack_1, ack => convTransposeD_CP_6059_elements(41)); -- 
    rr_6436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(41), ack => ptr_deref_2685_load_0_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Sample/word_access_start/$exit
      -- CP-element group 42: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Sample/word_access_start/word_0/$exit
      -- CP-element group 42: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Sample/word_access_start/word_0/ra
      -- 
    ra_6437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2685_load_0_ack_0, ack => convTransposeD_CP_6059_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	92 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	51 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Update/word_access_complete/$exit
      -- CP-element group 43: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Update/word_access_complete/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Update/word_access_complete/word_0/ca
      -- CP-element group 43: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Update/ptr_deref_2685_Merge/$entry
      -- CP-element group 43: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Update/ptr_deref_2685_Merge/$exit
      -- CP-element group 43: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Update/ptr_deref_2685_Merge/merge_req
      -- CP-element group 43: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Update/ptr_deref_2685_Merge/merge_ack
      -- 
    ca_6448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2685_load_0_ack_1, ack => convTransposeD_CP_6059_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	31 
    -- CP-element group 44: 	33 
    -- CP-element group 44: 	35 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2695_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2695_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2695_Sample/rr
      -- 
    rr_6461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(44), ack => type_cast_2695_inst_req_0); -- 
    convTransposeD_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(31) & convTransposeD_CP_6059_elements(33) & convTransposeD_CP_6059_elements(35);
      gj_convTransposeD_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2695_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2695_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2695_Sample/ra
      -- 
    ra_6462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2695_inst_ack_0, ack => convTransposeD_CP_6059_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	92 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (16) 
      -- CP-element group 46: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_index_scale_1/scale_rename_ack
      -- CP-element group 46: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_index_resized_1
      -- CP-element group 46: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_index_scale_1/scale_rename_req
      -- CP-element group 46: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_index_scale_1/$exit
      -- CP-element group 46: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_index_scale_1/$entry
      -- CP-element group 46: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_index_scaled_1
      -- CP-element group 46: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_final_index_sum_regn_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_index_computed_1
      -- CP-element group 46: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_index_resize_1/$entry
      -- CP-element group 46: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_final_index_sum_regn_Sample/req
      -- CP-element group 46: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_index_resize_1/index_resize_ack
      -- CP-element group 46: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_index_resize_1/index_resize_req
      -- CP-element group 46: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_index_resize_1/$exit
      -- CP-element group 46: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2695_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2695_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2695_Update/ca
      -- 
    ca_6467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2695_inst_ack_1, ack => convTransposeD_CP_6059_elements(46)); -- 
    req_6492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(46), ack => array_obj_ref_2701_index_offset_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	54 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_final_index_sum_regn_sample_complete
      -- CP-element group 47: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_final_index_sum_regn_Sample/ack
      -- CP-element group 47: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_final_index_sum_regn_Sample/$exit
      -- 
    ack_6493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2701_index_offset_ack_0, ack => convTransposeD_CP_6059_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	92 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (11) 
      -- CP-element group 48: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2702_request/$entry
      -- CP-element group 48: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2702_request/req
      -- CP-element group 48: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_root_address_calculated
      -- CP-element group 48: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_offset_calculated
      -- CP-element group 48: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_base_plus_offset/sum_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_base_plus_offset/sum_rename_req
      -- CP-element group 48: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_base_plus_offset/$exit
      -- CP-element group 48: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_base_plus_offset/$entry
      -- CP-element group 48: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_final_index_sum_regn_Update/ack
      -- CP-element group 48: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_final_index_sum_regn_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2702_sample_start_
      -- 
    ack_6498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2701_index_offset_ack_1, ack => convTransposeD_CP_6059_elements(48)); -- 
    req_6507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(48), ack => addr_of_2702_final_reg_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2702_request/$exit
      -- CP-element group 49: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2702_request/ack
      -- CP-element group 49: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2702_sample_completed_
      -- 
    ack_6508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2702_final_reg_ack_0, ack => convTransposeD_CP_6059_elements(49)); -- 
    -- CP-element group 50:  fork  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	92 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (19) 
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2702_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_base_addr_resize/base_resize_req
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_base_addr_resize/$entry
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_base_address_resized
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_base_addr_resize/$exit
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2702_complete/ack
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_base_addr_resize/base_resize_ack
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_base_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_word_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_word_addrgen/root_register_ack
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_word_addrgen/root_register_req
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_word_addrgen/$exit
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_word_addrgen/$entry
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_base_plus_offset/sum_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2702_update_completed_
      -- 
    ack_6513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2702_final_reg_ack_1, ack => convTransposeD_CP_6059_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	43 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Sample/word_access_start/word_0/rr
      -- CP-element group 51: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Sample/ptr_deref_2705_Split/split_ack
      -- CP-element group 51: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Sample/ptr_deref_2705_Split/split_req
      -- CP-element group 51: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Sample/ptr_deref_2705_Split/$exit
      -- CP-element group 51: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Sample/ptr_deref_2705_Split/$entry
      -- CP-element group 51: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Sample/$entry
      -- 
    rr_6551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(51), ack => ptr_deref_2705_store_0_req_0); -- 
    convTransposeD_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(43) & convTransposeD_CP_6059_elements(50);
      gj_convTransposeD_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Sample/word_access_start/word_0/ra
      -- CP-element group 52: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Sample/$exit
      -- 
    ra_6552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2705_store_0_ack_0, ack => convTransposeD_CP_6059_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	92 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Update/word_access_complete/word_0/ca
      -- CP-element group 53: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_update_completed_
      -- 
    ca_6563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2705_store_0_ack_1, ack => convTransposeD_CP_6059_elements(53)); -- 
    -- CP-element group 54:  branch  join  transition  place  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	38 
    -- CP-element group 54: 	47 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (10) 
      -- CP-element group 54: 	 branch_block_stmt_2429/if_stmt_2719_dead_link/$entry
      -- CP-element group 54: 	 branch_block_stmt_2429/if_stmt_2719_else_link/$entry
      -- CP-element group 54: 	 branch_block_stmt_2429/if_stmt_2719__entry__
      -- CP-element group 54: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718__exit__
      -- CP-element group 54: 	 branch_block_stmt_2429/R_cmp_2720_place
      -- CP-element group 54: 	 branch_block_stmt_2429/if_stmt_2719_eval_test/$entry
      -- CP-element group 54: 	 branch_block_stmt_2429/if_stmt_2719_eval_test/$exit
      -- CP-element group 54: 	 branch_block_stmt_2429/if_stmt_2719_eval_test/branch_req
      -- CP-element group 54: 	 branch_block_stmt_2429/if_stmt_2719_if_link/$entry
      -- CP-element group 54: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/$exit
      -- 
    branch_req_6571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(54), ack => if_stmt_2719_branch_req_0); -- 
    convTransposeD_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(38) & convTransposeD_CP_6059_elements(47) & convTransposeD_CP_6059_elements(53);
      gj_convTransposeD_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	101 
    -- CP-element group 55: 	102 
    -- CP-element group 55: 	104 
    -- CP-element group 55: 	105 
    -- CP-element group 55: 	107 
    -- CP-element group 55: 	108 
    -- CP-element group 55:  members (40) 
      -- CP-element group 55: 	 branch_block_stmt_2429/assign_stmt_2731/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138
      -- CP-element group 55: 	 branch_block_stmt_2429/assign_stmt_2731__exit__
      -- CP-element group 55: 	 branch_block_stmt_2429/assign_stmt_2731__entry__
      -- CP-element group 55: 	 branch_block_stmt_2429/whilex_xbody_ifx_xthen
      -- CP-element group 55: 	 branch_block_stmt_2429/merge_stmt_2725__exit__
      -- CP-element group 55: 	 branch_block_stmt_2429/assign_stmt_2731/$exit
      -- CP-element group 55: 	 branch_block_stmt_2429/merge_stmt_2725_PhiReqMerge
      -- CP-element group 55: 	 branch_block_stmt_2429/if_stmt_2719_if_link/$exit
      -- CP-element group 55: 	 branch_block_stmt_2429/if_stmt_2719_if_link/if_choice_transition
      -- CP-element group 55: 	 branch_block_stmt_2429/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 55: 	 branch_block_stmt_2429/merge_stmt_2725_PhiAck/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/merge_stmt_2725_PhiAck/$exit
      -- CP-element group 55: 	 branch_block_stmt_2429/merge_stmt_2725_PhiAck/dummy
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2781/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_sources/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_sources/type_cast_2784/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_sources/type_cast_2784/SplitProtocol/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_sources/type_cast_2784/SplitProtocol/Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_sources/type_cast_2784/SplitProtocol/Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_sources/type_cast_2784/SplitProtocol/Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_sources/type_cast_2784/SplitProtocol/Update/cr
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2788/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2791/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2791/SplitProtocol/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2791/SplitProtocol/Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2791/SplitProtocol/Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2791/SplitProtocol/Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2791/SplitProtocol/Update/cr
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2794/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2797/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2797/SplitProtocol/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2797/SplitProtocol/Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2797/SplitProtocol/Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2797/SplitProtocol/Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2797/SplitProtocol/Update/cr
      -- 
    if_choice_transition_6576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2719_branch_ack_1, ack => convTransposeD_CP_6059_elements(55)); -- 
    rr_6922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(55), ack => type_cast_2784_inst_req_0); -- 
    cr_6927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(55), ack => type_cast_2784_inst_req_1); -- 
    rr_6945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(55), ack => type_cast_2791_inst_req_0); -- 
    cr_6950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(55), ack => type_cast_2791_inst_req_1); -- 
    rr_6968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(55), ack => type_cast_2797_inst_req_0); -- 
    cr_6973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(55), ack => type_cast_2797_inst_req_1); -- 
    -- CP-element group 56:  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	58 
    -- CP-element group 56: 	60 
    -- CP-element group 56: 	62 
    -- CP-element group 56:  members (24) 
      -- CP-element group 56: 	 branch_block_stmt_2429/whilex_xbody_ifx_xelse
      -- CP-element group 56: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2751_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2751_update_start_
      -- CP-element group 56: 	 branch_block_stmt_2429/if_stmt_2719_else_link/else_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773__entry__
      -- CP-element group 56: 	 branch_block_stmt_2429/merge_stmt_2733__exit__
      -- CP-element group 56: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2767_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_2429/if_stmt_2719_else_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2767_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/$entry
      -- CP-element group 56: 	 branch_block_stmt_2429/merge_stmt_2733_PhiReqMerge
      -- CP-element group 56: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2751_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2742_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2767_update_start_
      -- CP-element group 56: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2742_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2742_Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2742_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2742_update_start_
      -- CP-element group 56: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2742_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_2429/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_2429/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_2429/merge_stmt_2733_PhiAck/$entry
      -- CP-element group 56: 	 branch_block_stmt_2429/merge_stmt_2733_PhiAck/$exit
      -- CP-element group 56: 	 branch_block_stmt_2429/merge_stmt_2733_PhiAck/dummy
      -- 
    else_choice_transition_6580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2719_branch_ack_0, ack => convTransposeD_CP_6059_elements(56)); -- 
    cr_6615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(56), ack => type_cast_2751_inst_req_1); -- 
    cr_6629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(56), ack => type_cast_2767_inst_req_1); -- 
    cr_6601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(56), ack => type_cast_2742_inst_req_1); -- 
    rr_6596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(56), ack => type_cast_2742_inst_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2742_Sample/ra
      -- CP-element group 57: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2742_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2742_sample_completed_
      -- 
    ra_6597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2742_inst_ack_0, ack => convTransposeD_CP_6059_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2742_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2751_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2751_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2751_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2742_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2742_update_completed_
      -- 
    ca_6602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2742_inst_ack_1, ack => convTransposeD_CP_6059_elements(58)); -- 
    rr_6610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(58), ack => type_cast_2751_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2751_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2751_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2751_Sample/ra
      -- 
    ra_6611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2751_inst_ack_0, ack => convTransposeD_CP_6059_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	56 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2751_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2767_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2767_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2751_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2767_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2751_Update/$exit
      -- 
    ca_6616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2751_inst_ack_1, ack => convTransposeD_CP_6059_elements(60)); -- 
    rr_6624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(60), ack => type_cast_2767_inst_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2767_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2767_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2767_sample_completed_
      -- 
    ra_6625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2767_inst_ack_0, ack => convTransposeD_CP_6059_elements(61)); -- 
    -- CP-element group 62:  branch  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	56 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (13) 
      -- CP-element group 62: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2767_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_2429/R_cmp127_2775_place
      -- CP-element group 62: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2767_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_2429/if_stmt_2774__entry__
      -- CP-element group 62: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773__exit__
      -- CP-element group 62: 	 branch_block_stmt_2429/if_stmt_2774_else_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_2429/if_stmt_2774_if_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_2429/if_stmt_2774_eval_test/branch_req
      -- CP-element group 62: 	 branch_block_stmt_2429/if_stmt_2774_eval_test/$exit
      -- CP-element group 62: 	 branch_block_stmt_2429/if_stmt_2774_eval_test/$entry
      -- CP-element group 62: 	 branch_block_stmt_2429/if_stmt_2774_dead_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/$exit
      -- CP-element group 62: 	 branch_block_stmt_2429/assign_stmt_2739_to_assign_stmt_2773/type_cast_2767_Update/$exit
      -- 
    ca_6630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2767_inst_ack_1, ack => convTransposeD_CP_6059_elements(62)); -- 
    branch_req_6638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(62), ack => if_stmt_2774_branch_req_0); -- 
    -- CP-element group 63:  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (15) 
      -- CP-element group 63: 	 branch_block_stmt_2429/ifx_xelse_whilex_xend
      -- CP-element group 63: 	 branch_block_stmt_2429/assign_stmt_2813__entry__
      -- CP-element group 63: 	 branch_block_stmt_2429/merge_stmt_2808__exit__
      -- CP-element group 63: 	 branch_block_stmt_2429/merge_stmt_2808_PhiReqMerge
      -- CP-element group 63: 	 branch_block_stmt_2429/assign_stmt_2813/WPIPE_Block3_done_2810_Sample/req
      -- CP-element group 63: 	 branch_block_stmt_2429/assign_stmt_2813/WPIPE_Block3_done_2810_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_2429/assign_stmt_2813/WPIPE_Block3_done_2810_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_2429/assign_stmt_2813/$entry
      -- CP-element group 63: 	 branch_block_stmt_2429/if_stmt_2774_if_link/if_choice_transition
      -- CP-element group 63: 	 branch_block_stmt_2429/if_stmt_2774_if_link/$exit
      -- CP-element group 63: 	 branch_block_stmt_2429/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 63: 	 branch_block_stmt_2429/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 63: 	 branch_block_stmt_2429/merge_stmt_2808_PhiAck/$entry
      -- CP-element group 63: 	 branch_block_stmt_2429/merge_stmt_2808_PhiAck/$exit
      -- CP-element group 63: 	 branch_block_stmt_2429/merge_stmt_2808_PhiAck/dummy
      -- 
    if_choice_transition_6643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2774_branch_ack_1, ack => convTransposeD_CP_6059_elements(63)); -- 
    req_6663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(63), ack => WPIPE_Block3_done_2810_inst_req_0); -- 
    -- CP-element group 64:  fork  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	93 
    -- CP-element group 64: 	94 
    -- CP-element group 64: 	95 
    -- CP-element group 64: 	97 
    -- CP-element group 64: 	98 
    -- CP-element group 64:  members (22) 
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138
      -- CP-element group 64: 	 branch_block_stmt_2429/if_stmt_2774_else_link/else_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_2429/if_stmt_2774_else_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2781/$entry
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_sources/$entry
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2788/$entry
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/$entry
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2793/$entry
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2793/SplitProtocol/$entry
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2793/SplitProtocol/Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2793/SplitProtocol/Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2793/SplitProtocol/Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2793/SplitProtocol/Update/cr
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2794/$entry
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/$entry
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2799/$entry
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2799/SplitProtocol/$entry
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2799/SplitProtocol/Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2799/SplitProtocol/Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2799/SplitProtocol/Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2799/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2774_branch_ack_0, ack => convTransposeD_CP_6059_elements(64)); -- 
    rr_6873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(64), ack => type_cast_2793_inst_req_0); -- 
    cr_6878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(64), ack => type_cast_2793_inst_req_1); -- 
    rr_6896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(64), ack => type_cast_2799_inst_req_0); -- 
    cr_6901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(64), ack => type_cast_2799_inst_req_1); -- 
    -- CP-element group 65:  transition  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (6) 
      -- CP-element group 65: 	 branch_block_stmt_2429/assign_stmt_2813/WPIPE_Block3_done_2810_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_2429/assign_stmt_2813/WPIPE_Block3_done_2810_Update/req
      -- CP-element group 65: 	 branch_block_stmt_2429/assign_stmt_2813/WPIPE_Block3_done_2810_Sample/ack
      -- CP-element group 65: 	 branch_block_stmt_2429/assign_stmt_2813/WPIPE_Block3_done_2810_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_2429/assign_stmt_2813/WPIPE_Block3_done_2810_update_start_
      -- CP-element group 65: 	 branch_block_stmt_2429/assign_stmt_2813/WPIPE_Block3_done_2810_sample_completed_
      -- 
    ack_6664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2810_inst_ack_0, ack => convTransposeD_CP_6059_elements(65)); -- 
    req_6668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(65), ack => WPIPE_Block3_done_2810_inst_req_1); -- 
    -- CP-element group 66:  transition  place  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (16) 
      -- CP-element group 66: 	 branch_block_stmt_2429/branch_block_stmt_2429__exit__
      -- CP-element group 66: 	 branch_block_stmt_2429/$exit
      -- CP-element group 66: 	 $exit
      -- CP-element group 66: 	 branch_block_stmt_2429/assign_stmt_2813/WPIPE_Block3_done_2810_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_2429/assign_stmt_2813__exit__
      -- CP-element group 66: 	 branch_block_stmt_2429/return__
      -- CP-element group 66: 	 branch_block_stmt_2429/merge_stmt_2815__exit__
      -- CP-element group 66: 	 branch_block_stmt_2429/assign_stmt_2813/WPIPE_Block3_done_2810_Update/ack
      -- CP-element group 66: 	 branch_block_stmt_2429/assign_stmt_2813/WPIPE_Block3_done_2810_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_2429/assign_stmt_2813/$exit
      -- CP-element group 66: 	 branch_block_stmt_2429/return___PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_2429/return___PhiReq/$exit
      -- CP-element group 66: 	 branch_block_stmt_2429/merge_stmt_2815_PhiReqMerge
      -- CP-element group 66: 	 branch_block_stmt_2429/merge_stmt_2815_PhiAck/$entry
      -- CP-element group 66: 	 branch_block_stmt_2429/merge_stmt_2815_PhiAck/$exit
      -- CP-element group 66: 	 branch_block_stmt_2429/merge_stmt_2815_PhiAck/dummy
      -- 
    ack_6669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_2810_inst_ack_1, ack => convTransposeD_CP_6059_elements(66)); -- 
    -- CP-element group 67:  transition  output  delay-element  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	29 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	73 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/$exit
      -- CP-element group 67: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2569_konst_delay_trans
      -- CP-element group 67: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_req
      -- CP-element group 67: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2563/$exit
      -- 
    phi_stmt_2563_req_6680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2563_req_6680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(67), ack => phi_stmt_2563_req_1); -- 
    -- Element group convTransposeD_CP_6059_elements(67) is a control-delay.
    cp_element_67_delay: control_delay_element  generic map(name => " 67_delay", delay_value => 1)  port map(req => convTransposeD_CP_6059_elements(29), ack => convTransposeD_CP_6059_elements(67), clk => clk, reset =>reset);
    -- CP-element group 68:  transition  output  delay-element  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	29 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	73 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_sources/type_cast_2576_konst_delay_trans
      -- CP-element group 68: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_req
      -- CP-element group 68: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2570/$exit
      -- CP-element group 68: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_sources/$exit
      -- 
    phi_stmt_2570_req_6688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2570_req_6688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(68), ack => phi_stmt_2570_req_1); -- 
    -- Element group convTransposeD_CP_6059_elements(68) is a control-delay.
    cp_element_68_delay: control_delay_element  generic map(name => " 68_delay", delay_value => 1)  port map(req => convTransposeD_CP_6059_elements(29), ack => convTransposeD_CP_6059_elements(68), clk => clk, reset =>reset);
    -- CP-element group 69:  transition  output  delay-element  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	29 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	73 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_sources/$exit
      -- CP-element group 69: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2577/$exit
      -- CP-element group 69: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_sources/type_cast_2583_konst_delay_trans
      -- CP-element group 69: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_req
      -- 
    phi_stmt_2577_req_6696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2577_req_6696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(69), ack => phi_stmt_2577_req_1); -- 
    -- Element group convTransposeD_CP_6059_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => convTransposeD_CP_6059_elements(29), ack => convTransposeD_CP_6059_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	29 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2587/SplitProtocol/Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2587/SplitProtocol/Sample/ra
      -- 
    ra_6713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2587_inst_ack_0, ack => convTransposeD_CP_6059_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	29 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2587/SplitProtocol/Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2587/SplitProtocol/Update/ca
      -- 
    ca_6718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2587_inst_ack_1, ack => convTransposeD_CP_6059_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (5) 
      -- CP-element group 72: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2584/$exit
      -- CP-element group 72: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/$exit
      -- CP-element group 72: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2587/$exit
      -- CP-element group 72: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2587/SplitProtocol/$exit
      -- CP-element group 72: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_req
      -- 
    phi_stmt_2584_req_6719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2584_req_6719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(72), ack => phi_stmt_2584_req_0); -- 
    convTransposeD_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(70) & convTransposeD_CP_6059_elements(71);
      gj_convTransposeD_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	67 
    -- CP-element group 73: 	68 
    -- CP-element group 73: 	69 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	87 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_2429/entry_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(67) & convTransposeD_CP_6059_elements(68) & convTransposeD_CP_6059_elements(69) & convTransposeD_CP_6059_elements(72);
      gj_convTransposeD_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	1 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Sample/ra
      -- 
    ra_6739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2566_inst_ack_0, ack => convTransposeD_CP_6059_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	1 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/Update/ca
      -- 
    ca_6744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2566_inst_ack_1, ack => convTransposeD_CP_6059_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	86 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2563/$exit
      -- CP-element group 76: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/$exit
      -- CP-element group 76: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_sources/type_cast_2566/SplitProtocol/$exit
      -- CP-element group 76: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2563/phi_stmt_2563_req
      -- 
    phi_stmt_2563_req_6745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2563_req_6745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(76), ack => phi_stmt_2563_req_0); -- 
    convTransposeD_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(74) & convTransposeD_CP_6059_elements(75);
      gj_convTransposeD_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	1 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_sources/type_cast_2573/SplitProtocol/Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_sources/type_cast_2573/SplitProtocol/Sample/ra
      -- 
    ra_6762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2573_inst_ack_0, ack => convTransposeD_CP_6059_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	1 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_sources/type_cast_2573/SplitProtocol/Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_sources/type_cast_2573/SplitProtocol/Update/ca
      -- 
    ca_6767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2573_inst_ack_1, ack => convTransposeD_CP_6059_elements(78)); -- 
    -- CP-element group 79:  join  transition  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	86 
    -- CP-element group 79:  members (5) 
      -- CP-element group 79: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2570/$exit
      -- CP-element group 79: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_sources/$exit
      -- CP-element group 79: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_sources/type_cast_2573/$exit
      -- CP-element group 79: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_sources/type_cast_2573/SplitProtocol/$exit
      -- CP-element group 79: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2570/phi_stmt_2570_req
      -- 
    phi_stmt_2570_req_6768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2570_req_6768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(79), ack => phi_stmt_2570_req_0); -- 
    convTransposeD_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(77) & convTransposeD_CP_6059_elements(78);
      gj_convTransposeD_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	1 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_sources/type_cast_2580/SplitProtocol/Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_sources/type_cast_2580/SplitProtocol/Sample/ra
      -- 
    ra_6785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2580_inst_ack_0, ack => convTransposeD_CP_6059_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	1 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_sources/type_cast_2580/SplitProtocol/Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_sources/type_cast_2580/SplitProtocol/Update/ca
      -- 
    ca_6790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2580_inst_ack_1, ack => convTransposeD_CP_6059_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	86 
    -- CP-element group 82:  members (5) 
      -- CP-element group 82: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2577/$exit
      -- CP-element group 82: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_sources/$exit
      -- CP-element group 82: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_sources/type_cast_2580/$exit
      -- CP-element group 82: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_sources/type_cast_2580/SplitProtocol/$exit
      -- CP-element group 82: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2577/phi_stmt_2577_req
      -- 
    phi_stmt_2577_req_6791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2577_req_6791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(82), ack => phi_stmt_2577_req_0); -- 
    convTransposeD_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(80) & convTransposeD_CP_6059_elements(81);
      gj_convTransposeD_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	1 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2589/SplitProtocol/Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2589/SplitProtocol/Sample/ra
      -- 
    ra_6808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2589_inst_ack_0, ack => convTransposeD_CP_6059_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	1 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2589/SplitProtocol/Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2589/SplitProtocol/Update/ca
      -- 
    ca_6813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2589_inst_ack_1, ack => convTransposeD_CP_6059_elements(84)); -- 
    -- CP-element group 85:  join  transition  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2584/$exit
      -- CP-element group 85: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/$exit
      -- CP-element group 85: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2589/$exit
      -- CP-element group 85: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_sources/type_cast_2589/SplitProtocol/$exit
      -- CP-element group 85: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/phi_stmt_2584/phi_stmt_2584_req
      -- 
    phi_stmt_2584_req_6814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2584_req_6814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(85), ack => phi_stmt_2584_req_1); -- 
    convTransposeD_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(83) & convTransposeD_CP_6059_elements(84);
      gj_convTransposeD_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  join  transition  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	76 
    -- CP-element group 86: 	79 
    -- CP-element group 86: 	82 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_2429/ifx_xend138_whilex_xbody_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(76) & convTransposeD_CP_6059_elements(79) & convTransposeD_CP_6059_elements(82) & convTransposeD_CP_6059_elements(85);
      gj_convTransposeD_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  merge  fork  transition  place  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	73 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	89 
    -- CP-element group 87: 	90 
    -- CP-element group 87: 	91 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2429/merge_stmt_2562_PhiReqMerge
      -- CP-element group 87: 	 branch_block_stmt_2429/merge_stmt_2562_PhiAck/$entry
      -- 
    convTransposeD_CP_6059_elements(87) <= OrReduce(convTransposeD_CP_6059_elements(73) & convTransposeD_CP_6059_elements(86));
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	92 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_2429/merge_stmt_2562_PhiAck/phi_stmt_2563_ack
      -- 
    phi_stmt_2563_ack_6819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2563_ack_0, ack => convTransposeD_CP_6059_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	92 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_2429/merge_stmt_2562_PhiAck/phi_stmt_2570_ack
      -- 
    phi_stmt_2570_ack_6820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2570_ack_0, ack => convTransposeD_CP_6059_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_2429/merge_stmt_2562_PhiAck/phi_stmt_2577_ack
      -- 
    phi_stmt_2577_ack_6821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2577_ack_0, ack => convTransposeD_CP_6059_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	87 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_2429/merge_stmt_2562_PhiAck/phi_stmt_2584_ack
      -- 
    phi_stmt_2584_ack_6822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2584_ack_0, ack => convTransposeD_CP_6059_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  place  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	88 
    -- CP-element group 92: 	89 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	30 
    -- CP-element group 92: 	31 
    -- CP-element group 92: 	32 
    -- CP-element group 92: 	33 
    -- CP-element group 92: 	34 
    -- CP-element group 92: 	35 
    -- CP-element group 92: 	36 
    -- CP-element group 92: 	37 
    -- CP-element group 92: 	39 
    -- CP-element group 92: 	41 
    -- CP-element group 92: 	43 
    -- CP-element group 92: 	46 
    -- CP-element group 92: 	48 
    -- CP-element group 92: 	50 
    -- CP-element group 92: 	53 
    -- CP-element group 92:  members (53) 
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2702_complete/req
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/merge_stmt_2562__exit__
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718__entry__
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Update/word_access_complete/word_0/cr
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_final_index_sum_regn_update_start
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2702_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Update/word_access_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2705_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_final_index_sum_regn_Update/req
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2701_final_index_sum_regn_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2604_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2604_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2604_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2604_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2604_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2604_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2618_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2618_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2618_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2618_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2618_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2618_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2632_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2632_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2632_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2632_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2632_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2632_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2674_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2674_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2674_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2674_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2674_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2674_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2681_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_final_index_sum_regn_update_start
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_final_index_sum_regn_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/array_obj_ref_2680_final_index_sum_regn_Update/req
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2681_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2681_complete/req
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Update/word_access_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/ptr_deref_2685_Update/word_access_complete/word_0/cr
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2695_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2695_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/type_cast_2695_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2429/assign_stmt_2596_to_assign_stmt_2718/addr_of_2702_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2429/merge_stmt_2562_PhiAck/$exit
      -- 
    req_6512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(92), ack => addr_of_2702_final_reg_req_1); -- 
    cr_6562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(92), ack => ptr_deref_2705_store_0_req_1); -- 
    req_6497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(92), ack => array_obj_ref_2701_index_offset_req_1); -- 
    rr_6309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(92), ack => type_cast_2604_inst_req_0); -- 
    cr_6314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(92), ack => type_cast_2604_inst_req_1); -- 
    rr_6323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(92), ack => type_cast_2618_inst_req_0); -- 
    cr_6328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(92), ack => type_cast_2618_inst_req_1); -- 
    rr_6337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(92), ack => type_cast_2632_inst_req_0); -- 
    cr_6342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(92), ack => type_cast_2632_inst_req_1); -- 
    rr_6351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(92), ack => type_cast_2674_inst_req_0); -- 
    cr_6356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(92), ack => type_cast_2674_inst_req_1); -- 
    req_6387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(92), ack => array_obj_ref_2680_index_offset_req_1); -- 
    req_6402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(92), ack => addr_of_2681_final_reg_req_1); -- 
    cr_6447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(92), ack => ptr_deref_2685_load_0_req_1); -- 
    cr_6466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(92), ack => type_cast_2695_inst_req_1); -- 
    convTransposeD_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(88) & convTransposeD_CP_6059_elements(89) & convTransposeD_CP_6059_elements(90) & convTransposeD_CP_6059_elements(91);
      gj_convTransposeD_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  output  delay-element  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	64 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	100 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2781/$exit
      -- CP-element group 93: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_sources/$exit
      -- CP-element group 93: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_sources/type_cast_2787_konst_delay_trans
      -- CP-element group 93: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_req
      -- 
    phi_stmt_2781_req_6857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2781_req_6857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(93), ack => phi_stmt_2781_req_1); -- 
    -- Element group convTransposeD_CP_6059_elements(93) is a control-delay.
    cp_element_93_delay: control_delay_element  generic map(name => " 93_delay", delay_value => 1)  port map(req => convTransposeD_CP_6059_elements(64), ack => convTransposeD_CP_6059_elements(93), clk => clk, reset =>reset);
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	64 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2793/SplitProtocol/Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2793/SplitProtocol/Sample/ra
      -- 
    ra_6874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2793_inst_ack_0, ack => convTransposeD_CP_6059_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	64 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2793/SplitProtocol/Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2793/SplitProtocol/Update/ca
      -- 
    ca_6879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2793_inst_ack_1, ack => convTransposeD_CP_6059_elements(95)); -- 
    -- CP-element group 96:  join  transition  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	100 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2788/$exit
      -- CP-element group 96: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/$exit
      -- CP-element group 96: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2793/$exit
      -- CP-element group 96: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2793/SplitProtocol/$exit
      -- CP-element group 96: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_req
      -- 
    phi_stmt_2788_req_6880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2788_req_6880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(96), ack => phi_stmt_2788_req_1); -- 
    convTransposeD_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(94) & convTransposeD_CP_6059_elements(95);
      gj_convTransposeD_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	64 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2799/SplitProtocol/Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2799/SplitProtocol/Sample/ra
      -- 
    ra_6897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2799_inst_ack_0, ack => convTransposeD_CP_6059_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	64 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2799/SplitProtocol/Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2799/SplitProtocol/Update/ca
      -- 
    ca_6902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2799_inst_ack_1, ack => convTransposeD_CP_6059_elements(98)); -- 
    -- CP-element group 99:  join  transition  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2794/$exit
      -- CP-element group 99: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/$exit
      -- CP-element group 99: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2799/$exit
      -- CP-element group 99: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2799/SplitProtocol/$exit
      -- CP-element group 99: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_req
      -- 
    phi_stmt_2794_req_6903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2794_req_6903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(99), ack => phi_stmt_2794_req_1); -- 
    convTransposeD_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(97) & convTransposeD_CP_6059_elements(98);
      gj_convTransposeD_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  join  transition  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	93 
    -- CP-element group 100: 	96 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	111 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_2429/ifx_xelse_ifx_xend138_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(93) & convTransposeD_CP_6059_elements(96) & convTransposeD_CP_6059_elements(99);
      gj_convTransposeD_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	55 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_sources/type_cast_2784/SplitProtocol/Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_sources/type_cast_2784/SplitProtocol/Sample/ra
      -- 
    ra_6923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2784_inst_ack_0, ack => convTransposeD_CP_6059_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	55 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_sources/type_cast_2784/SplitProtocol/Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_sources/type_cast_2784/SplitProtocol/Update/ca
      -- 
    ca_6928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2784_inst_ack_1, ack => convTransposeD_CP_6059_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	110 
    -- CP-element group 103:  members (5) 
      -- CP-element group 103: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2781/$exit
      -- CP-element group 103: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_sources/$exit
      -- CP-element group 103: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_sources/type_cast_2784/$exit
      -- CP-element group 103: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_sources/type_cast_2784/SplitProtocol/$exit
      -- CP-element group 103: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2781/phi_stmt_2781_req
      -- 
    phi_stmt_2781_req_6929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2781_req_6929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(103), ack => phi_stmt_2781_req_0); -- 
    convTransposeD_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(101) & convTransposeD_CP_6059_elements(102);
      gj_convTransposeD_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	55 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2791/SplitProtocol/Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2791/SplitProtocol/Sample/ra
      -- 
    ra_6946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2791_inst_ack_0, ack => convTransposeD_CP_6059_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	55 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2791/SplitProtocol/Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2791/SplitProtocol/Update/ca
      -- 
    ca_6951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2791_inst_ack_1, ack => convTransposeD_CP_6059_elements(105)); -- 
    -- CP-element group 106:  join  transition  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	110 
    -- CP-element group 106:  members (5) 
      -- CP-element group 106: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2788/$exit
      -- CP-element group 106: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/$exit
      -- CP-element group 106: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2791/$exit
      -- CP-element group 106: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_sources/type_cast_2791/SplitProtocol/$exit
      -- CP-element group 106: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2788/phi_stmt_2788_req
      -- 
    phi_stmt_2788_req_6952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2788_req_6952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(106), ack => phi_stmt_2788_req_0); -- 
    convTransposeD_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(104) & convTransposeD_CP_6059_elements(105);
      gj_convTransposeD_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	55 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2797/SplitProtocol/Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2797/SplitProtocol/Sample/ra
      -- 
    ra_6969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2797_inst_ack_0, ack => convTransposeD_CP_6059_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	55 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2797/SplitProtocol/Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2797/SplitProtocol/Update/ca
      -- 
    ca_6974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2797_inst_ack_1, ack => convTransposeD_CP_6059_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2794/$exit
      -- CP-element group 109: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/$exit
      -- CP-element group 109: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2797/$exit
      -- CP-element group 109: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_sources/type_cast_2797/SplitProtocol/$exit
      -- CP-element group 109: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/phi_stmt_2794/phi_stmt_2794_req
      -- 
    phi_stmt_2794_req_6975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2794_req_6975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_6059_elements(109), ack => phi_stmt_2794_req_0); -- 
    convTransposeD_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(107) & convTransposeD_CP_6059_elements(108);
      gj_convTransposeD_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  transition  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	103 
    -- CP-element group 110: 	106 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_2429/ifx_xthen_ifx_xend138_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(103) & convTransposeD_CP_6059_elements(106) & convTransposeD_CP_6059_elements(109);
      gj_convTransposeD_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  merge  fork  transition  place  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	100 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	113 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_2429/merge_stmt_2780_PhiReqMerge
      -- CP-element group 111: 	 branch_block_stmt_2429/merge_stmt_2780_PhiAck/$entry
      -- 
    convTransposeD_CP_6059_elements(111) <= OrReduce(convTransposeD_CP_6059_elements(100) & convTransposeD_CP_6059_elements(110));
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	115 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2429/merge_stmt_2780_PhiAck/phi_stmt_2781_ack
      -- 
    phi_stmt_2781_ack_6980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2781_ack_0, ack => convTransposeD_CP_6059_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_2429/merge_stmt_2780_PhiAck/phi_stmt_2788_ack
      -- 
    phi_stmt_2788_ack_6981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2788_ack_0, ack => convTransposeD_CP_6059_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_2429/merge_stmt_2780_PhiAck/phi_stmt_2794_ack
      -- 
    phi_stmt_2794_ack_6982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2794_ack_0, ack => convTransposeD_CP_6059_elements(114)); -- 
    -- CP-element group 115:  join  transition  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	112 
    -- CP-element group 115: 	113 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	1 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_2429/merge_stmt_2780_PhiAck/$exit
      -- 
    convTransposeD_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convTransposeD_CP_6059_elements(112) & convTransposeD_CP_6059_elements(113) & convTransposeD_CP_6059_elements(114);
      gj_convTransposeD_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_6059_elements(115), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_idxprom97_2700_resized : std_logic_vector(13 downto 0);
    signal R_idxprom97_2700_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2679_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2679_scaled : std_logic_vector(13 downto 0);
    signal add102_2713 : std_logic_vector(31 downto 0);
    signal add109_2731 : std_logic_vector(15 downto 0);
    signal add56_2514 : std_logic_vector(31 downto 0);
    signal add69_2525 : std_logic_vector(31 downto 0);
    signal add88_2655 : std_logic_vector(31 downto 0);
    signal add90_2665 : std_logic_vector(31 downto 0);
    signal add_2498 : std_logic_vector(31 downto 0);
    signal add_src_0x_x0_2601 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2680_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2680_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2680_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2680_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2680_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2680_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2701_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2701_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2701_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2701_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2701_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2701_root_address : std_logic_vector(13 downto 0);
    signal arrayidx93_2682 : std_logic_vector(31 downto 0);
    signal arrayidx98_2703 : std_logic_vector(31 downto 0);
    signal call10_2444 : std_logic_vector(31 downto 0);
    signal call13_2447 : std_logic_vector(31 downto 0);
    signal call16_2450 : std_logic_vector(31 downto 0);
    signal call19_2453 : std_logic_vector(31 downto 0);
    signal call1_2435 : std_logic_vector(31 downto 0);
    signal call21_2456 : std_logic_vector(31 downto 0);
    signal call23_2459 : std_logic_vector(31 downto 0);
    signal call24_2462 : std_logic_vector(31 downto 0);
    signal call27_2465 : std_logic_vector(31 downto 0);
    signal call30_2468 : std_logic_vector(31 downto 0);
    signal call4_2438 : std_logic_vector(31 downto 0);
    signal call7_2441 : std_logic_vector(31 downto 0);
    signal call_2432 : std_logic_vector(31 downto 0);
    signal cmp117_2748 : std_logic_vector(0 downto 0);
    signal cmp127_2773 : std_logic_vector(0 downto 0);
    signal cmp_2718 : std_logic_vector(0 downto 0);
    signal conv105_2548 : std_logic_vector(31 downto 0);
    signal conv113_2743 : std_logic_vector(31 downto 0);
    signal conv116_2554 : std_logic_vector(31 downto 0);
    signal conv123_2768 : std_logic_vector(31 downto 0);
    signal conv126_2560 : std_logic_vector(31 downto 0);
    signal conv34_2475 : std_logic_vector(31 downto 0);
    signal conv37_2487 : std_logic_vector(31 downto 0);
    signal conv39_2502 : std_logic_vector(15 downto 0);
    signal conv50_2605 : std_logic_vector(31 downto 0);
    signal conv52_2508 : std_logic_vector(31 downto 0);
    signal conv62_2619 : std_logic_vector(31 downto 0);
    signal conv76_2633 : std_logic_vector(31 downto 0);
    signal conv79_2536 : std_logic_vector(31 downto 0);
    signal conv81_2639 : std_logic_vector(31 downto 0);
    signal conv84_2542 : std_logic_vector(31 downto 0);
    signal conv86_2645 : std_logic_vector(31 downto 0);
    signal idxprom97_2696 : std_logic_vector(63 downto 0);
    signal idxprom_2675 : std_logic_vector(63 downto 0);
    signal inc121_2752 : std_logic_vector(15 downto 0);
    signal inc121x_xinput_dim0x_x2_2757 : std_logic_vector(15 downto 0);
    signal inc_2739 : std_logic_vector(15 downto 0);
    signal indvar_2563 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_2806 : std_logic_vector(31 downto 0);
    signal input_dim0x_x1x_xph_2794 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2_2584 : std_logic_vector(15 downto 0);
    signal input_dim1x_x0x_xph_2788 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1_2577 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2764 : std_logic_vector(15 downto 0);
    signal input_dim2x_x0x_xph_2781 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2570 : std_logic_vector(15 downto 0);
    signal mul65_2624 : std_logic_vector(31 downto 0);
    signal mul87_2650 : std_logic_vector(31 downto 0);
    signal mul89_2660 : std_logic_vector(31 downto 0);
    signal mul_2610 : std_logic_vector(31 downto 0);
    signal ptr_deref_2685_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2685_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2685_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2685_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2685_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2705_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2705_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2705_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2705_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2705_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2705_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr141_2481 : std_logic_vector(31 downto 0);
    signal shr38142_2493 : std_logic_vector(31 downto 0);
    signal shr92_2671 : std_logic_vector(31 downto 0);
    signal shr96_2692 : std_logic_vector(31 downto 0);
    signal sub59_2615 : std_logic_vector(31 downto 0);
    signal sub72_2530 : std_logic_vector(31 downto 0);
    signal sub73_2629 : std_logic_vector(31 downto 0);
    signal sub_2519 : std_logic_vector(31 downto 0);
    signal tmp1_2596 : std_logic_vector(31 downto 0);
    signal tmp94_2686 : std_logic_vector(63 downto 0);
    signal type_cast_2473_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2479_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2485_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2491_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2506_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2512_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2523_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2534_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2540_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2546_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2552_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2558_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2566_wire : std_logic_vector(31 downto 0);
    signal type_cast_2569_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2573_wire : std_logic_vector(15 downto 0);
    signal type_cast_2576_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2580_wire : std_logic_vector(15 downto 0);
    signal type_cast_2583_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2587_wire : std_logic_vector(15 downto 0);
    signal type_cast_2589_wire : std_logic_vector(15 downto 0);
    signal type_cast_2594_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2637_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2643_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2669_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2690_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2711_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2729_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2737_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2761_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2784_wire : std_logic_vector(15 downto 0);
    signal type_cast_2787_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2791_wire : std_logic_vector(15 downto 0);
    signal type_cast_2793_wire : std_logic_vector(15 downto 0);
    signal type_cast_2797_wire : std_logic_vector(15 downto 0);
    signal type_cast_2799_wire : std_logic_vector(15 downto 0);
    signal type_cast_2804_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2812_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_2680_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2680_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2680_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2680_resized_base_address <= "00000000000000";
    array_obj_ref_2701_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2701_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2701_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2701_resized_base_address <= "00000000000000";
    ptr_deref_2685_word_offset_0 <= "00000000000000";
    ptr_deref_2705_word_offset_0 <= "00000000000000";
    type_cast_2473_wire_constant <= "00000000000000000000000000000010";
    type_cast_2479_wire_constant <= "00000000000000000011111111111111";
    type_cast_2485_wire_constant <= "00000000000000000000000000000001";
    type_cast_2491_wire_constant <= "00000000000000000111111111111111";
    type_cast_2506_wire_constant <= "00000000000000001111111111111111";
    type_cast_2512_wire_constant <= "00000000000000001111111111111111";
    type_cast_2523_wire_constant <= "00000000000000001111111111111111";
    type_cast_2534_wire_constant <= "00000000000000001111111111111111";
    type_cast_2540_wire_constant <= "00000000000000001111111111111111";
    type_cast_2546_wire_constant <= "00000000000000001111111111111111";
    type_cast_2552_wire_constant <= "00000000000000001111111111111111";
    type_cast_2558_wire_constant <= "00000000000000001111111111111111";
    type_cast_2569_wire_constant <= "00000000000000000000000000000000";
    type_cast_2576_wire_constant <= "0000000000000000";
    type_cast_2583_wire_constant <= "0000000000000000";
    type_cast_2594_wire_constant <= "00000000000000000000000000000100";
    type_cast_2637_wire_constant <= "00000000000000001111111111111111";
    type_cast_2643_wire_constant <= "00000000000000001111111111111111";
    type_cast_2669_wire_constant <= "00000000000000000000000000000010";
    type_cast_2690_wire_constant <= "00000000000000000000000000000010";
    type_cast_2711_wire_constant <= "00000000000000000000000000000100";
    type_cast_2729_wire_constant <= "0000000000000100";
    type_cast_2737_wire_constant <= "0000000000000001";
    type_cast_2761_wire_constant <= "0000000000000000";
    type_cast_2787_wire_constant <= "0000000000000000";
    type_cast_2804_wire_constant <= "00000000000000000000000000000001";
    type_cast_2812_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_2563: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2566_wire & type_cast_2569_wire_constant;
      req <= phi_stmt_2563_req_0 & phi_stmt_2563_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2563",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2563_ack_0,
          idata => idata,
          odata => indvar_2563,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2563
    phi_stmt_2570: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2573_wire & type_cast_2576_wire_constant;
      req <= phi_stmt_2570_req_0 & phi_stmt_2570_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2570",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2570_ack_0,
          idata => idata,
          odata => input_dim2x_x1_2570,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2570
    phi_stmt_2577: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2580_wire & type_cast_2583_wire_constant;
      req <= phi_stmt_2577_req_0 & phi_stmt_2577_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2577",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2577_ack_0,
          idata => idata,
          odata => input_dim1x_x1_2577,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2577
    phi_stmt_2584: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2587_wire & type_cast_2589_wire;
      req <= phi_stmt_2584_req_0 & phi_stmt_2584_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2584",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2584_ack_0,
          idata => idata,
          odata => input_dim0x_x2_2584,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2584
    phi_stmt_2781: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2784_wire & type_cast_2787_wire_constant;
      req <= phi_stmt_2781_req_0 & phi_stmt_2781_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2781",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2781_ack_0,
          idata => idata,
          odata => input_dim2x_x0x_xph_2781,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2781
    phi_stmt_2788: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2791_wire & type_cast_2793_wire;
      req <= phi_stmt_2788_req_0 & phi_stmt_2788_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2788",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2788_ack_0,
          idata => idata,
          odata => input_dim1x_x0x_xph_2788,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2788
    phi_stmt_2794: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2797_wire & type_cast_2799_wire;
      req <= phi_stmt_2794_req_0 & phi_stmt_2794_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2794",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2794_ack_0,
          idata => idata,
          odata => input_dim0x_x1x_xph_2794,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2794
    -- flow-through select operator MUX_2763_inst
    input_dim1x_x2_2764 <= type_cast_2761_wire_constant when (cmp117_2748(0) /=  '0') else inc_2739;
    addr_of_2681_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2681_final_reg_req_0;
      addr_of_2681_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2681_final_reg_req_1;
      addr_of_2681_final_reg_ack_1<= rack(0);
      addr_of_2681_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2681_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2680_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx93_2682,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2702_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2702_final_reg_req_0;
      addr_of_2702_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2702_final_reg_req_1;
      addr_of_2702_final_reg_ack_1<= rack(0);
      addr_of_2702_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2702_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2701_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx98_2703,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2501_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2501_inst_req_0;
      type_cast_2501_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2501_inst_req_1;
      type_cast_2501_inst_ack_1<= rack(0);
      type_cast_2501_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2501_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_2498,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_2502,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2566_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2566_inst_req_0;
      type_cast_2566_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2566_inst_req_1;
      type_cast_2566_inst_ack_1<= rack(0);
      type_cast_2566_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2566_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2806,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2566_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2573_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2573_inst_req_0;
      type_cast_2573_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2573_inst_req_1;
      type_cast_2573_inst_ack_1<= rack(0);
      type_cast_2573_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2573_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x0x_xph_2781,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2573_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2580_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2580_inst_req_0;
      type_cast_2580_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2580_inst_req_1;
      type_cast_2580_inst_ack_1<= rack(0);
      type_cast_2580_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2580_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x0x_xph_2788,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2580_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2587_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2587_inst_req_0;
      type_cast_2587_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2587_inst_req_1;
      type_cast_2587_inst_ack_1<= rack(0);
      type_cast_2587_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2587_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv39_2502,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2587_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2589_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2589_inst_req_0;
      type_cast_2589_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2589_inst_req_1;
      type_cast_2589_inst_ack_1<= rack(0);
      type_cast_2589_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2589_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x1x_xph_2794,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2589_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2604_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2604_inst_req_0;
      type_cast_2604_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2604_inst_req_1;
      type_cast_2604_inst_ack_1<= rack(0);
      type_cast_2604_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2604_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2584,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv50_2605,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2618_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2618_inst_req_0;
      type_cast_2618_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2618_inst_req_1;
      type_cast_2618_inst_ack_1<= rack(0);
      type_cast_2618_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2618_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2577,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_2619,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2632_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2632_inst_req_0;
      type_cast_2632_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2632_inst_req_1;
      type_cast_2632_inst_ack_1<= rack(0);
      type_cast_2632_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2632_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2570,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv76_2633,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2674_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2674_inst_req_0;
      type_cast_2674_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2674_inst_req_1;
      type_cast_2674_inst_ack_1<= rack(0);
      type_cast_2674_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2674_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr92_2671,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2675,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2695_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2695_inst_req_0;
      type_cast_2695_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2695_inst_req_1;
      type_cast_2695_inst_ack_1<= rack(0);
      type_cast_2695_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2695_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr96_2692,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom97_2696,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2742_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2742_inst_req_0;
      type_cast_2742_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2742_inst_req_1;
      type_cast_2742_inst_ack_1<= rack(0);
      type_cast_2742_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2742_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_2739,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_2743,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2751_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2751_inst_req_0;
      type_cast_2751_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2751_inst_req_1;
      type_cast_2751_inst_ack_1<= rack(0);
      type_cast_2751_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2751_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp117_2748,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc121_2752,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2767_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2767_inst_req_0;
      type_cast_2767_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2767_inst_req_1;
      type_cast_2767_inst_ack_1<= rack(0);
      type_cast_2767_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2767_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc121x_xinput_dim0x_x2_2757,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv123_2768,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2784_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2784_inst_req_0;
      type_cast_2784_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2784_inst_req_1;
      type_cast_2784_inst_ack_1<= rack(0);
      type_cast_2784_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2784_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add109_2731,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2784_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2791_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2791_inst_req_0;
      type_cast_2791_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2791_inst_req_1;
      type_cast_2791_inst_ack_1<= rack(0);
      type_cast_2791_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2791_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x1_2577,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2791_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2793_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2793_inst_req_0;
      type_cast_2793_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2793_inst_req_1;
      type_cast_2793_inst_ack_1<= rack(0);
      type_cast_2793_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2793_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2764,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2793_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2797_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2797_inst_req_0;
      type_cast_2797_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2797_inst_req_1;
      type_cast_2797_inst_ack_1<= rack(0);
      type_cast_2797_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2797_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2_2584,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2797_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2799_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2799_inst_req_0;
      type_cast_2799_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2799_inst_req_1;
      type_cast_2799_inst_ack_1<= rack(0);
      type_cast_2799_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2799_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc121x_xinput_dim0x_x2_2757,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2799_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_2680_index_1_rename
    process(R_idxprom_2679_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2679_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2679_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2680_index_1_resize
    process(idxprom_2675) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2675;
      ov := iv(13 downto 0);
      R_idxprom_2679_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2680_root_address_inst
    process(array_obj_ref_2680_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2680_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2680_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2701_index_1_rename
    process(R_idxprom97_2700_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom97_2700_resized;
      ov(13 downto 0) := iv;
      R_idxprom97_2700_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2701_index_1_resize
    process(idxprom97_2696) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom97_2696;
      ov := iv(13 downto 0);
      R_idxprom97_2700_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2701_root_address_inst
    process(array_obj_ref_2701_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2701_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2701_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2685_addr_0
    process(ptr_deref_2685_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2685_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2685_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2685_base_resize
    process(arrayidx93_2682) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx93_2682;
      ov := iv(13 downto 0);
      ptr_deref_2685_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2685_gather_scatter
    process(ptr_deref_2685_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2685_data_0;
      ov(63 downto 0) := iv;
      tmp94_2686 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2685_root_address_inst
    process(ptr_deref_2685_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2685_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2685_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2705_addr_0
    process(ptr_deref_2705_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2705_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2705_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2705_base_resize
    process(arrayidx98_2703) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx98_2703;
      ov := iv(13 downto 0);
      ptr_deref_2705_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2705_gather_scatter
    process(tmp94_2686) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp94_2686;
      ov(63 downto 0) := iv;
      ptr_deref_2705_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2705_root_address_inst
    process(ptr_deref_2705_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2705_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2705_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2719_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2718;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2719_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2719_branch_req_0,
          ack0 => if_stmt_2719_branch_ack_0,
          ack1 => if_stmt_2719_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2774_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp127_2773;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2774_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2774_branch_req_0,
          ack0 => if_stmt_2774_branch_ack_0,
          ack1 => if_stmt_2774_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2730_inst
    process(input_dim2x_x1_2570) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim2x_x1_2570, type_cast_2729_wire_constant, tmp_var);
      add109_2731 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2738_inst
    process(input_dim1x_x1_2577) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1_2577, type_cast_2737_wire_constant, tmp_var);
      inc_2739 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2756_inst
    process(inc121_2752, input_dim0x_x2_2584) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc121_2752, input_dim0x_x2_2584, tmp_var);
      inc121x_xinput_dim0x_x2_2757 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2497_inst
    process(shr141_2481, shr38142_2493) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr141_2481, shr38142_2493, tmp_var);
      add_2498 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2513_inst
    process(call10_2444) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call10_2444, type_cast_2512_wire_constant, tmp_var);
      add56_2514 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2524_inst
    process(call13_2447) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call13_2447, type_cast_2523_wire_constant, tmp_var);
      add69_2525 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2600_inst
    process(call23_2459, tmp1_2596) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(call23_2459, tmp1_2596, tmp_var);
      add_src_0x_x0_2601 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2614_inst
    process(sub_2519, mul_2610) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub_2519, mul_2610, tmp_var);
      sub59_2615 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2628_inst
    process(sub72_2530, mul65_2624) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub72_2530, mul65_2624, tmp_var);
      sub73_2629 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2654_inst
    process(mul87_2650, conv81_2639) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul87_2650, conv81_2639, tmp_var);
      add88_2655 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2664_inst
    process(mul89_2660, conv76_2633) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul89_2660, conv76_2633, tmp_var);
      add90_2665 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2712_inst
    process(conv76_2633) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv76_2633, type_cast_2711_wire_constant, tmp_var);
      add102_2713 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2805_inst
    process(indvar_2563) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2563, type_cast_2804_wire_constant, tmp_var);
      indvarx_xnext_2806 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2480_inst
    process(conv34_2475) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv34_2475, type_cast_2479_wire_constant, tmp_var);
      shr141_2481 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2492_inst
    process(conv37_2487) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv37_2487, type_cast_2491_wire_constant, tmp_var);
      shr38142_2493 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2507_inst
    process(call19_2453) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call19_2453, type_cast_2506_wire_constant, tmp_var);
      conv52_2508 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2535_inst
    process(call30_2468) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call30_2468, type_cast_2534_wire_constant, tmp_var);
      conv79_2536 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2541_inst
    process(call27_2465) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call27_2465, type_cast_2540_wire_constant, tmp_var);
      conv84_2542 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2547_inst
    process(call4_2438) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call4_2438, type_cast_2546_wire_constant, tmp_var);
      conv105_2548 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2553_inst
    process(call1_2435) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call1_2435, type_cast_2552_wire_constant, tmp_var);
      conv116_2554 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2559_inst
    process(call_2432) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(call_2432, type_cast_2558_wire_constant, tmp_var);
      conv126_2560 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2638_inst
    process(sub73_2629) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(sub73_2629, type_cast_2637_wire_constant, tmp_var);
      conv81_2639 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_2644_inst
    process(sub59_2615) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(sub59_2615, type_cast_2643_wire_constant, tmp_var);
      conv86_2645 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2747_inst
    process(conv113_2743, conv116_2554) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv113_2743, conv116_2554, tmp_var);
      cmp117_2748 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2772_inst
    process(conv123_2768, conv126_2560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv123_2768, conv126_2560, tmp_var);
      cmp127_2773 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2474_inst
    process(call_2432) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2432, type_cast_2473_wire_constant, tmp_var);
      conv34_2475 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2486_inst
    process(call_2432) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(call_2432, type_cast_2485_wire_constant, tmp_var);
      conv37_2487 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2670_inst
    process(add_src_0x_x0_2601) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add_src_0x_x0_2601, type_cast_2669_wire_constant, tmp_var);
      shr92_2671 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2691_inst
    process(add90_2665) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add90_2665, type_cast_2690_wire_constant, tmp_var);
      shr96_2692 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2595_inst
    process(indvar_2563) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2563, type_cast_2594_wire_constant, tmp_var);
      tmp1_2596 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2609_inst
    process(conv50_2605, conv52_2508) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv50_2605, conv52_2508, tmp_var);
      mul_2610 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2623_inst
    process(conv62_2619, conv52_2508) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv62_2619, conv52_2508, tmp_var);
      mul65_2624 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2649_inst
    process(conv86_2645, conv84_2542) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv86_2645, conv84_2542, tmp_var);
      mul87_2650 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2659_inst
    process(add88_2655, conv79_2536) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add88_2655, conv79_2536, tmp_var);
      mul89_2660 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2518_inst
    process(add56_2514, call21_2456) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add56_2514, call21_2456, tmp_var);
      sub_2519 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2529_inst
    process(add69_2525, call21_2456) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add69_2525, call21_2456, tmp_var);
      sub72_2530 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2717_inst
    process(add102_2713, conv105_2548) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add102_2713, conv105_2548, tmp_var);
      cmp_2718 <= tmp_var; --
    end process;
    -- shared split operator group (37) : array_obj_ref_2680_index_offset 
    ApIntAdd_group_37: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2679_scaled;
      array_obj_ref_2680_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2680_index_offset_req_0;
      array_obj_ref_2680_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2680_index_offset_req_1;
      array_obj_ref_2680_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_37_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_37_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_37",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : array_obj_ref_2701_index_offset 
    ApIntAdd_group_38: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom97_2700_scaled;
      array_obj_ref_2701_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2701_index_offset_req_0;
      array_obj_ref_2701_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2701_index_offset_req_1;
      array_obj_ref_2701_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_38_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_38_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_38",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared load operator group (0) : ptr_deref_2685_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2685_load_0_req_0;
      ptr_deref_2685_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2685_load_0_req_1;
      ptr_deref_2685_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2685_word_address_0;
      ptr_deref_2685_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_2705_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2705_store_0_req_0;
      ptr_deref_2705_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2705_store_0_req_1;
      ptr_deref_2705_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2705_word_address_0;
      data_in <= ptr_deref_2705_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2431_inst RPIPE_Block3_start_2434_inst RPIPE_Block3_start_2437_inst RPIPE_Block3_start_2440_inst RPIPE_Block3_start_2443_inst RPIPE_Block3_start_2446_inst RPIPE_Block3_start_2449_inst RPIPE_Block3_start_2452_inst RPIPE_Block3_start_2455_inst RPIPE_Block3_start_2458_inst RPIPE_Block3_start_2461_inst RPIPE_Block3_start_2464_inst RPIPE_Block3_start_2467_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(415 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 12 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 12 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 12 downto 0);
      signal guard_vector : std_logic_vector( 12 downto 0);
      constant outBUFs : IntegerArray(12 downto 0) := (12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(12 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false);
      constant guardBuffering: IntegerArray(12 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2);
      -- 
    begin -- 
      reqL_unguarded(12) <= RPIPE_Block3_start_2431_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Block3_start_2434_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Block3_start_2437_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Block3_start_2440_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Block3_start_2443_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Block3_start_2446_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Block3_start_2449_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block3_start_2452_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block3_start_2455_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block3_start_2458_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block3_start_2461_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block3_start_2464_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block3_start_2467_inst_req_0;
      RPIPE_Block3_start_2431_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Block3_start_2434_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Block3_start_2437_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Block3_start_2440_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Block3_start_2443_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Block3_start_2446_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Block3_start_2449_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block3_start_2452_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block3_start_2455_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block3_start_2458_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block3_start_2461_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block3_start_2464_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block3_start_2467_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(12) <= RPIPE_Block3_start_2431_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Block3_start_2434_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Block3_start_2437_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Block3_start_2440_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Block3_start_2443_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Block3_start_2446_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Block3_start_2449_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block3_start_2452_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block3_start_2455_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block3_start_2458_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block3_start_2461_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block3_start_2464_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block3_start_2467_inst_req_1;
      RPIPE_Block3_start_2431_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Block3_start_2434_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Block3_start_2437_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Block3_start_2440_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Block3_start_2443_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Block3_start_2446_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Block3_start_2449_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block3_start_2452_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block3_start_2455_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block3_start_2458_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block3_start_2461_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block3_start_2464_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block3_start_2467_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      call_2432 <= data_out(415 downto 384);
      call1_2435 <= data_out(383 downto 352);
      call4_2438 <= data_out(351 downto 320);
      call7_2441 <= data_out(319 downto 288);
      call10_2444 <= data_out(287 downto 256);
      call13_2447 <= data_out(255 downto 224);
      call16_2450 <= data_out(223 downto 192);
      call19_2453 <= data_out(191 downto 160);
      call21_2456 <= data_out(159 downto 128);
      call23_2459 <= data_out(127 downto 96);
      call24_2462 <= data_out(95 downto 64);
      call27_2465 <= data_out(63 downto 32);
      call30_2468 <= data_out(31 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 13, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 32,  num_reqs => 13,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_2810_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_2810_inst_req_0;
      WPIPE_Block3_done_2810_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_2810_inst_req_1;
      WPIPE_Block3_done_2810_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_2812_wire_constant;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_28_load_0_req_0 : boolean;
  signal LOAD_count_28_load_0_ack_0 : boolean;
  signal LOAD_count_28_load_0_req_1 : boolean;
  signal LOAD_count_28_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_29/$entry
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_sample_start_
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_update_start_
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_29/LOAD_count_28_Sample/$entry
      -- 
    rr_21_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_21_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_28_load_0_req_0); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => LOAD_count_28_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_sample_completed_
      -- CP-element group 1: 	 assign_stmt_29/LOAD_count_28_Sample/$exit
      -- 
    ra_22_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_28_load_0_ack_0, ack => timer_CP_0_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/$entry
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_29/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_update_completed_
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_29/LOAD_count_28_Update/LOAD_count_28_Merge/merge_ack
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_28_load_0_ack_1, ack => timer_CP_0_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_28_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_28_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_28_word_address_0 <= "0";
    -- equivalence LOAD_count_28_gather_scatter
    process(LOAD_count_28_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_28_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_28_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_28_load_0_req_0;
      LOAD_count_28_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_28_load_0_req_1;
      LOAD_count_28_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_28_word_address_0;
      LOAD_count_28_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(4 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(31 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(31 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(31 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(31 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(31 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(31 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(31 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(31 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(31 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(31 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(31 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(31 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(31 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(31 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(31 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(31 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(31 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(31 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(31 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(31 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(31 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(31 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(31 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(31 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(31 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(31 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(31 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(31 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(18 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(0 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(10 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(0 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(4 downto 4),
      memory_space_3_sr_ack => memory_space_3_sr_ack(4 downto 4),
      memory_space_3_sr_addr => memory_space_3_sr_addr(69 downto 56),
      memory_space_3_sr_data => memory_space_3_sr_data(319 downto 256),
      memory_space_3_sr_tag => memory_space_3_sr_tag(94 downto 76),
      memory_space_3_sc_req => memory_space_3_sc_req(4 downto 4),
      memory_space_3_sc_ack => memory_space_3_sc_ack(4 downto 4),
      memory_space_3_sc_tag => memory_space_3_sc_tag(4 downto 4),
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(31 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(31 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(31 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(31 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(31 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(31 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(31 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(31 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(55 downto 42),
      memory_space_1_lr_tag => memory_space_1_lr_tag(75 downto 57),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(255 downto 192),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 3),
      memory_space_3_sr_req => memory_space_3_sr_req(3 downto 3),
      memory_space_3_sr_ack => memory_space_3_sr_ack(3 downto 3),
      memory_space_3_sr_addr => memory_space_3_sr_addr(55 downto 42),
      memory_space_3_sr_data => memory_space_3_sr_data(255 downto 192),
      memory_space_3_sr_tag => memory_space_3_sr_tag(75 downto 57),
      memory_space_3_sc_req => memory_space_3_sc_req(3 downto 3),
      memory_space_3_sc_ack => memory_space_3_sc_ack(3 downto 3),
      memory_space_3_sc_tag => memory_space_3_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(31 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(31 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(41 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(56 downto 38),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(191 downto 128),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 2),
      memory_space_3_sr_req => memory_space_3_sr_req(2 downto 2),
      memory_space_3_sr_ack => memory_space_3_sr_ack(2 downto 2),
      memory_space_3_sr_addr => memory_space_3_sr_addr(41 downto 28),
      memory_space_3_sr_data => memory_space_3_sr_data(191 downto 128),
      memory_space_3_sr_tag => memory_space_3_sr_tag(56 downto 38),
      memory_space_3_sc_req => memory_space_3_sc_req(2 downto 2),
      memory_space_3_sc_ack => memory_space_3_sc_ack(2 downto 2),
      memory_space_3_sc_tag => memory_space_3_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(31 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(31 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(13 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(18 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(0 downto 0),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(31 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(31 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(37 downto 19),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(127 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 1),
      memory_space_3_sr_req => memory_space_3_sr_req(1 downto 1),
      memory_space_3_sr_ack => memory_space_3_sr_ack(1 downto 1),
      memory_space_3_sr_addr => memory_space_3_sr_addr(27 downto 14),
      memory_space_3_sr_data => memory_space_3_sr_data(127 downto 64),
      memory_space_3_sr_tag => memory_space_3_sr_tag(37 downto 19),
      memory_space_3_sc_req => memory_space_3_sc_req(1 downto 1),
      memory_space_3_sc_ack => memory_space_3_sc_ack(1 downto 1),
      memory_space_3_sc_tag => memory_space_3_sc_tag(1 downto 1),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(31 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(31 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(0 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  dummyROM_memory_space_0: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_2: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
